module hann(input logic [11:0] n, output logic [23:0] coeff);
    always_comb begin
        case(n)
            12'd0: coeff = 24'd0;
            12'd1: coeff = 24'd9;
            12'd2: coeff = 24'd39;
            12'd3: coeff = 24'd88;
            12'd4: coeff = 24'd157;
            12'd5: coeff = 24'd246;
            12'd6: coeff = 24'd355;
            12'd7: coeff = 24'd483;
            12'd8: coeff = 24'd631;
            12'd9: coeff = 24'd799;
            12'd10: coeff = 24'd987;
            12'd11: coeff = 24'd1194;
            12'd12: coeff = 24'd1421;
            12'd13: coeff = 24'd1668;
            12'd14: coeff = 24'd1935;
            12'd15: coeff = 24'd2221;
            12'd16: coeff = 24'd2527;
            12'd17: coeff = 24'd2853;
            12'd18: coeff = 24'd3199;
            12'd19: coeff = 24'd3564;
            12'd20: coeff = 24'd3949;
            12'd21: coeff = 24'd4354;
            12'd22: coeff = 24'd4778;
            12'd23: coeff = 24'd5223;
            12'd24: coeff = 24'd5687;
            12'd25: coeff = 24'd6170;
            12'd26: coeff = 24'd6674;
            12'd27: coeff = 24'd7197;
            12'd28: coeff = 24'd7740;
            12'd29: coeff = 24'd8303;
            12'd30: coeff = 24'd8885;
            12'd31: coeff = 24'd9487;
            12'd32: coeff = 24'd10109;
            12'd33: coeff = 24'd10750;
            12'd34: coeff = 24'd11412;
            12'd35: coeff = 24'd12093;
            12'd36: coeff = 24'd12794;
            12'd37: coeff = 24'd13514;
            12'd38: coeff = 24'd14254;
            12'd39: coeff = 24'd15014;
            12'd40: coeff = 24'd15794;
            12'd41: coeff = 24'd16593;
            12'd42: coeff = 24'd17412;
            12'd43: coeff = 24'd18251;
            12'd44: coeff = 24'd19109;
            12'd45: coeff = 24'd19987;
            12'd46: coeff = 24'd20885;
            12'd47: coeff = 24'd21803;
            12'd48: coeff = 24'd22740;
            12'd49: coeff = 24'd23697;
            12'd50: coeff = 24'd24673;
            12'd51: coeff = 24'd25670;
            12'd52: coeff = 24'd26686;
            12'd53: coeff = 24'd27721;
            12'd54: coeff = 24'd28777;
            12'd55: coeff = 24'd29852;
            12'd56: coeff = 24'd30947;
            12'd57: coeff = 24'd32061;
            12'd58: coeff = 24'd33195;
            12'd59: coeff = 24'd34349;
            12'd60: coeff = 24'd35522;
            12'd61: coeff = 24'd36715;
            12'd62: coeff = 24'd37928;
            12'd63: coeff = 24'd39161;
            12'd64: coeff = 24'd40413;
            12'd65: coeff = 24'd41684;
            12'd66: coeff = 24'd42976;
            12'd67: coeff = 24'd44287;
            12'd68: coeff = 24'd45617;
            12'd69: coeff = 24'd46968;
            12'd70: coeff = 24'd48338;
            12'd71: coeff = 24'd49727;
            12'd72: coeff = 24'd51136;
            12'd73: coeff = 24'd52565;
            12'd74: coeff = 24'd54014;
            12'd75: coeff = 24'd55482;
            12'd76: coeff = 24'd56970;
            12'd77: coeff = 24'd58477;
            12'd78: coeff = 24'd60004;
            12'd79: coeff = 24'd61550;
            12'd80: coeff = 24'd63117;
            12'd81: coeff = 24'd64702;
            12'd82: coeff = 24'd66308;
            12'd83: coeff = 24'd67933;
            12'd84: coeff = 24'd69577;
            12'd85: coeff = 24'd71241;
            12'd86: coeff = 24'd72925;
            12'd87: coeff = 24'd74628;
            12'd88: coeff = 24'd76351;
            12'd89: coeff = 24'd78093;
            12'd90: coeff = 24'd79855;
            12'd91: coeff = 24'd81637;
            12'd92: coeff = 24'd83438;
            12'd93: coeff = 24'd85259;
            12'd94: coeff = 24'd87099;
            12'd95: coeff = 24'd88959;
            12'd96: coeff = 24'd90838;
            12'd97: coeff = 24'd92737;
            12'd98: coeff = 24'd94655;
            12'd99: coeff = 24'd96593;
            12'd100: coeff = 24'd98550;
            12'd101: coeff = 24'd100527;
            12'd102: coeff = 24'd102523;
            12'd103: coeff = 24'd104539;
            12'd104: coeff = 24'd106575;
            12'd105: coeff = 24'd108630;
            12'd106: coeff = 24'd110704;
            12'd107: coeff = 24'd112798;
            12'd108: coeff = 24'd114911;
            12'd109: coeff = 24'd117044;
            12'd110: coeff = 24'd119197;
            12'd111: coeff = 24'd121368;
            12'd112: coeff = 24'd123560;
            12'd113: coeff = 24'd125770;
            12'd114: coeff = 24'd128001;
            12'd115: coeff = 24'd130250;
            12'd116: coeff = 24'd132519;
            12'd117: coeff = 24'd134808;
            12'd118: coeff = 24'd137116;
            12'd119: coeff = 24'd139443;
            12'd120: coeff = 24'd141790;
            12'd121: coeff = 24'd144156;
            12'd122: coeff = 24'd146542;
            12'd123: coeff = 24'd148947;
            12'd124: coeff = 24'd151371;
            12'd125: coeff = 24'd153815;
            12'd126: coeff = 24'd156278;
            12'd127: coeff = 24'd158761;
            12'd128: coeff = 24'd161263;
            12'd129: coeff = 24'd163784;
            12'd130: coeff = 24'd166325;
            12'd131: coeff = 24'd168885;
            12'd132: coeff = 24'd171464;
            12'd133: coeff = 24'd174063;
            12'd134: coeff = 24'd176681;
            12'd135: coeff = 24'd179318;
            12'd136: coeff = 24'd181975;
            12'd137: coeff = 24'd184651;
            12'd138: coeff = 24'd187347;
            12'd139: coeff = 24'd190061;
            12'd140: coeff = 24'd192795;
            12'd141: coeff = 24'd195548;
            12'd142: coeff = 24'd198321;
            12'd143: coeff = 24'd201113;
            12'd144: coeff = 24'd203924;
            12'd145: coeff = 24'd206754;
            12'd146: coeff = 24'd209604;
            12'd147: coeff = 24'd212473;
            12'd148: coeff = 24'd215361;
            12'd149: coeff = 24'd218268;
            12'd150: coeff = 24'd221195;
            12'd151: coeff = 24'd224141;
            12'd152: coeff = 24'd227106;
            12'd153: coeff = 24'd230090;
            12'd154: coeff = 24'd233094;
            12'd155: coeff = 24'd236117;
            12'd156: coeff = 24'd239158;
            12'd157: coeff = 24'd242219;
            12'd158: coeff = 24'd245300;
            12'd159: coeff = 24'd248399;
            12'd160: coeff = 24'd251518;
            12'd161: coeff = 24'd254655;
            12'd162: coeff = 24'd257812;
            12'd163: coeff = 24'd260988;
            12'd164: coeff = 24'd264184;
            12'd165: coeff = 24'd267398;
            12'd166: coeff = 24'd270631;
            12'd167: coeff = 24'd273884;
            12'd168: coeff = 24'd277156;
            12'd169: coeff = 24'd280446;
            12'd170: coeff = 24'd283756;
            12'd171: coeff = 24'd287085;
            12'd172: coeff = 24'd290433;
            12'd173: coeff = 24'd293800;
            12'd174: coeff = 24'd297186;
            12'd175: coeff = 24'd300591;
            12'd176: coeff = 24'd304015;
            12'd177: coeff = 24'd307459;
            12'd178: coeff = 24'd310921;
            12'd179: coeff = 24'd314402;
            12'd180: coeff = 24'd317902;
            12'd181: coeff = 24'd321422;
            12'd182: coeff = 24'd324960;
            12'd183: coeff = 24'd328517;
            12'd184: coeff = 24'd332093;
            12'd185: coeff = 24'd335689;
            12'd186: coeff = 24'd339303;
            12'd187: coeff = 24'd342936;
            12'd188: coeff = 24'd346588;
            12'd189: coeff = 24'd350259;
            12'd190: coeff = 24'd353949;
            12'd191: coeff = 24'd357658;
            12'd192: coeff = 24'd361385;
            12'd193: coeff = 24'd365132;
            12'd194: coeff = 24'd368897;
            12'd195: coeff = 24'd372682;
            12'd196: coeff = 24'd376485;
            12'd197: coeff = 24'd380307;
            12'd198: coeff = 24'd384148;
            12'd199: coeff = 24'd388008;
            12'd200: coeff = 24'd391887;
            12'd201: coeff = 24'd395784;
            12'd202: coeff = 24'd399700;
            12'd203: coeff = 24'd403636;
            12'd204: coeff = 24'd407589;
            12'd205: coeff = 24'd411562;
            12'd206: coeff = 24'd415554;
            12'd207: coeff = 24'd419564;
            12'd208: coeff = 24'd423593;
            12'd209: coeff = 24'd427641;
            12'd210: coeff = 24'd431707;
            12'd211: coeff = 24'd435792;
            12'd212: coeff = 24'd439896;
            12'd213: coeff = 24'd444019;
            12'd214: coeff = 24'd448160;
            12'd215: coeff = 24'd452320;
            12'd216: coeff = 24'd456499;
            12'd217: coeff = 24'd460697;
            12'd218: coeff = 24'd464913;
            12'd219: coeff = 24'd469147;
            12'd220: coeff = 24'd473401;
            12'd221: coeff = 24'd477673;
            12'd222: coeff = 24'd481963;
            12'd223: coeff = 24'd486273;
            12'd224: coeff = 24'd490601;
            12'd225: coeff = 24'd494947;
            12'd226: coeff = 24'd499312;
            12'd227: coeff = 24'd503696;
            12'd228: coeff = 24'd508098;
            12'd229: coeff = 24'd512519;
            12'd230: coeff = 24'd516958;
            12'd231: coeff = 24'd521416;
            12'd232: coeff = 24'd525892;
            12'd233: coeff = 24'd530387;
            12'd234: coeff = 24'd534900;
            12'd235: coeff = 24'd539432;
            12'd236: coeff = 24'd543982;
            12'd237: coeff = 24'd548551;
            12'd238: coeff = 24'd553138;
            12'd239: coeff = 24'd557744;
            12'd240: coeff = 24'd562368;
            12'd241: coeff = 24'd567011;
            12'd242: coeff = 24'd571672;
            12'd243: coeff = 24'd576351;
            12'd244: coeff = 24'd581049;
            12'd245: coeff = 24'd585765;
            12'd246: coeff = 24'd590499;
            12'd247: coeff = 24'd595252;
            12'd248: coeff = 24'd600023;
            12'd249: coeff = 24'd604813;
            12'd250: coeff = 24'd609621;
            12'd251: coeff = 24'd614447;
            12'd252: coeff = 24'd619291;
            12'd253: coeff = 24'd624154;
            12'd254: coeff = 24'd629035;
            12'd255: coeff = 24'd633935;
            12'd256: coeff = 24'd638852;
            12'd257: coeff = 24'd643788;
            12'd258: coeff = 24'd648742;
            12'd259: coeff = 24'd653714;
            12'd260: coeff = 24'd658705;
            12'd261: coeff = 24'd663713;
            12'd262: coeff = 24'd668740;
            12'd263: coeff = 24'd673785;
            12'd264: coeff = 24'd678849;
            12'd265: coeff = 24'd683930;
            12'd266: coeff = 24'd689029;
            12'd267: coeff = 24'd694147;
            12'd268: coeff = 24'd699283;
            12'd269: coeff = 24'd704437;
            12'd270: coeff = 24'd709609;
            12'd271: coeff = 24'd714799;
            12'd272: coeff = 24'd720007;
            12'd273: coeff = 24'd725233;
            12'd274: coeff = 24'd730477;
            12'd275: coeff = 24'd735739;
            12'd276: coeff = 24'd741019;
            12'd277: coeff = 24'd746318;
            12'd278: coeff = 24'd751634;
            12'd279: coeff = 24'd756968;
            12'd280: coeff = 24'd762320;
            12'd281: coeff = 24'd767690;
            12'd282: coeff = 24'd773078;
            12'd283: coeff = 24'd778484;
            12'd284: coeff = 24'd783908;
            12'd285: coeff = 24'd789350;
            12'd286: coeff = 24'd794810;
            12'd287: coeff = 24'd800287;
            12'd288: coeff = 24'd805783;
            12'd289: coeff = 24'd811296;
            12'd290: coeff = 24'd816827;
            12'd291: coeff = 24'd822376;
            12'd292: coeff = 24'd827943;
            12'd293: coeff = 24'd833527;
            12'd294: coeff = 24'd839130;
            12'd295: coeff = 24'd844750;
            12'd296: coeff = 24'd850388;
            12'd297: coeff = 24'd856043;
            12'd298: coeff = 24'd861717;
            12'd299: coeff = 24'd867408;
            12'd300: coeff = 24'd873117;
            12'd301: coeff = 24'd878843;
            12'd302: coeff = 24'd884587;
            12'd303: coeff = 24'd890349;
            12'd304: coeff = 24'd896129;
            12'd305: coeff = 24'd901926;
            12'd306: coeff = 24'd907740;
            12'd307: coeff = 24'd913573;
            12'd308: coeff = 24'd919423;
            12'd309: coeff = 24'd925290;
            12'd310: coeff = 24'd931175;
            12'd311: coeff = 24'd937078;
            12'd312: coeff = 24'd942998;
            12'd313: coeff = 24'd948936;
            12'd314: coeff = 24'd954891;
            12'd315: coeff = 24'd960864;
            12'd316: coeff = 24'd966854;
            12'd317: coeff = 24'd972862;
            12'd318: coeff = 24'd978887;
            12'd319: coeff = 24'd984930;
            12'd320: coeff = 24'd990990;
            12'd321: coeff = 24'd997067;
            12'd322: coeff = 24'd1003162;
            12'd323: coeff = 24'd1009274;
            12'd324: coeff = 24'd1015404;
            12'd325: coeff = 24'd1021551;
            12'd326: coeff = 24'd1027715;
            12'd327: coeff = 24'd1033897;
            12'd328: coeff = 24'd1040096;
            12'd329: coeff = 24'd1046312;
            12'd330: coeff = 24'd1052546;
            12'd331: coeff = 24'd1058797;
            12'd332: coeff = 24'd1065065;
            12'd333: coeff = 24'd1071350;
            12'd334: coeff = 24'd1077653;
            12'd335: coeff = 24'd1083972;
            12'd336: coeff = 24'd1090309;
            12'd337: coeff = 24'd1096663;
            12'd338: coeff = 24'd1103035;
            12'd339: coeff = 24'd1109423;
            12'd340: coeff = 24'd1115829;
            12'd341: coeff = 24'd1122252;
            12'd342: coeff = 24'd1128691;
            12'd343: coeff = 24'd1135148;
            12'd344: coeff = 24'd1141622;
            12'd345: coeff = 24'd1148113;
            12'd346: coeff = 24'd1154621;
            12'd347: coeff = 24'd1161147;
            12'd348: coeff = 24'd1167689;
            12'd349: coeff = 24'd1174248;
            12'd350: coeff = 24'd1180824;
            12'd351: coeff = 24'd1187417;
            12'd352: coeff = 24'd1194027;
            12'd353: coeff = 24'd1200654;
            12'd354: coeff = 24'd1207298;
            12'd355: coeff = 24'd1213959;
            12'd356: coeff = 24'd1220637;
            12'd357: coeff = 24'd1227331;
            12'd358: coeff = 24'd1234043;
            12'd359: coeff = 24'd1240771;
            12'd360: coeff = 24'd1247516;
            12'd361: coeff = 24'd1254278;
            12'd362: coeff = 24'd1261057;
            12'd363: coeff = 24'd1267852;
            12'd364: coeff = 24'd1274664;
            12'd365: coeff = 24'd1281493;
            12'd366: coeff = 24'd1288339;
            12'd367: coeff = 24'd1295202;
            12'd368: coeff = 24'd1302081;
            12'd369: coeff = 24'd1308977;
            12'd370: coeff = 24'd1315889;
            12'd371: coeff = 24'd1322818;
            12'd372: coeff = 24'd1329764;
            12'd373: coeff = 24'd1336727;
            12'd374: coeff = 24'd1343706;
            12'd375: coeff = 24'd1350701;
            12'd376: coeff = 24'd1357713;
            12'd377: coeff = 24'd1364742;
            12'd378: coeff = 24'd1371787;
            12'd379: coeff = 24'd1378849;
            12'd380: coeff = 24'd1385927;
            12'd381: coeff = 24'd1393022;
            12'd382: coeff = 24'd1400133;
            12'd383: coeff = 24'd1407261;
            12'd384: coeff = 24'd1414405;
            12'd385: coeff = 24'd1421566;
            12'd386: coeff = 24'd1428743;
            12'd387: coeff = 24'd1435936;
            12'd388: coeff = 24'd1443146;
            12'd389: coeff = 24'd1450372;
            12'd390: coeff = 24'd1457614;
            12'd391: coeff = 24'd1464873;
            12'd392: coeff = 24'd1472148;
            12'd393: coeff = 24'd1479439;
            12'd394: coeff = 24'd1486747;
            12'd395: coeff = 24'd1494071;
            12'd396: coeff = 24'd1501411;
            12'd397: coeff = 24'd1508767;
            12'd398: coeff = 24'd1516139;
            12'd399: coeff = 24'd1523528;
            12'd400: coeff = 24'd1530933;
            12'd401: coeff = 24'd1538354;
            12'd402: coeff = 24'd1545791;
            12'd403: coeff = 24'd1553244;
            12'd404: coeff = 24'd1560713;
            12'd405: coeff = 24'd1568199;
            12'd406: coeff = 24'd1575700;
            12'd407: coeff = 24'd1583217;
            12'd408: coeff = 24'd1590751;
            12'd409: coeff = 24'd1598300;
            12'd410: coeff = 24'd1605866;
            12'd411: coeff = 24'd1613447;
            12'd412: coeff = 24'd1621045;
            12'd413: coeff = 24'd1628658;
            12'd414: coeff = 24'd1636287;
            12'd415: coeff = 24'd1643932;
            12'd416: coeff = 24'd1651593;
            12'd417: coeff = 24'd1659270;
            12'd418: coeff = 24'd1666963;
            12'd419: coeff = 24'd1674671;
            12'd420: coeff = 24'd1682396;
            12'd421: coeff = 24'd1690136;
            12'd422: coeff = 24'd1697892;
            12'd423: coeff = 24'd1705663;
            12'd424: coeff = 24'd1713451;
            12'd425: coeff = 24'd1721254;
            12'd426: coeff = 24'd1729072;
            12'd427: coeff = 24'd1736907;
            12'd428: coeff = 24'd1744757;
            12'd429: coeff = 24'd1752623;
            12'd430: coeff = 24'd1760504;
            12'd431: coeff = 24'd1768401;
            12'd432: coeff = 24'd1776314;
            12'd433: coeff = 24'd1784242;
            12'd434: coeff = 24'd1792185;
            12'd435: coeff = 24'd1800145;
            12'd436: coeff = 24'd1808119;
            12'd437: coeff = 24'd1816110;
            12'd438: coeff = 24'd1824115;
            12'd439: coeff = 24'd1832136;
            12'd440: coeff = 24'd1840173;
            12'd441: coeff = 24'd1848225;
            12'd442: coeff = 24'd1856292;
            12'd443: coeff = 24'd1864375;
            12'd444: coeff = 24'd1872473;
            12'd445: coeff = 24'd1880587;
            12'd446: coeff = 24'd1888716;
            12'd447: coeff = 24'd1896860;
            12'd448: coeff = 24'd1905019;
            12'd449: coeff = 24'd1913194;
            12'd450: coeff = 24'd1921384;
            12'd451: coeff = 24'd1929589;
            12'd452: coeff = 24'd1937809;
            12'd453: coeff = 24'd1946044;
            12'd454: coeff = 24'd1954295;
            12'd455: coeff = 24'd1962561;
            12'd456: coeff = 24'd1970842;
            12'd457: coeff = 24'd1979138;
            12'd458: coeff = 24'd1987449;
            12'd459: coeff = 24'd1995775;
            12'd460: coeff = 24'd2004117;
            12'd461: coeff = 24'd2012473;
            12'd462: coeff = 24'd2020844;
            12'd463: coeff = 24'd2029230;
            12'd464: coeff = 24'd2037632;
            12'd465: coeff = 24'd2046048;
            12'd466: coeff = 24'd2054479;
            12'd467: coeff = 24'd2062925;
            12'd468: coeff = 24'd2071386;
            12'd469: coeff = 24'd2079862;
            12'd470: coeff = 24'd2088353;
            12'd471: coeff = 24'd2096858;
            12'd472: coeff = 24'd2105379;
            12'd473: coeff = 24'd2113914;
            12'd474: coeff = 24'd2122464;
            12'd475: coeff = 24'd2131028;
            12'd476: coeff = 24'd2139608;
            12'd477: coeff = 24'd2148202;
            12'd478: coeff = 24'd2156810;
            12'd479: coeff = 24'd2165434;
            12'd480: coeff = 24'd2174072;
            12'd481: coeff = 24'd2182725;
            12'd482: coeff = 24'd2191392;
            12'd483: coeff = 24'd2200074;
            12'd484: coeff = 24'd2208771;
            12'd485: coeff = 24'd2217482;
            12'd486: coeff = 24'd2226207;
            12'd487: coeff = 24'd2234947;
            12'd488: coeff = 24'd2243702;
            12'd489: coeff = 24'd2252471;
            12'd490: coeff = 24'd2261254;
            12'd491: coeff = 24'd2270052;
            12'd492: coeff = 24'd2278865;
            12'd493: coeff = 24'd2287691;
            12'd494: coeff = 24'd2296532;
            12'd495: coeff = 24'd2305388;
            12'd496: coeff = 24'd2314257;
            12'd497: coeff = 24'd2323141;
            12'd498: coeff = 24'd2332040;
            12'd499: coeff = 24'd2340952;
            12'd500: coeff = 24'd2349879;
            12'd501: coeff = 24'd2358820;
            12'd502: coeff = 24'd2367775;
            12'd503: coeff = 24'd2376745;
            12'd504: coeff = 24'd2385728;
            12'd505: coeff = 24'd2394726;
            12'd506: coeff = 24'd2403738;
            12'd507: coeff = 24'd2412764;
            12'd508: coeff = 24'd2421804;
            12'd509: coeff = 24'd2430858;
            12'd510: coeff = 24'd2439926;
            12'd511: coeff = 24'd2449008;
            12'd512: coeff = 24'd2458104;
            12'd513: coeff = 24'd2467214;
            12'd514: coeff = 24'd2476338;
            12'd515: coeff = 24'd2485475;
            12'd516: coeff = 24'd2494627;
            12'd517: coeff = 24'd2503793;
            12'd518: coeff = 24'd2512972;
            12'd519: coeff = 24'd2522165;
            12'd520: coeff = 24'd2531373;
            12'd521: coeff = 24'd2540593;
            12'd522: coeff = 24'd2549828;
            12'd523: coeff = 24'd2559076;
            12'd524: coeff = 24'd2568339;
            12'd525: coeff = 24'd2577614;
            12'd526: coeff = 24'd2586904;
            12'd527: coeff = 24'd2596207;
            12'd528: coeff = 24'd2605524;
            12'd529: coeff = 24'd2614854;
            12'd530: coeff = 24'd2624198;
            12'd531: coeff = 24'd2633556;
            12'd532: coeff = 24'd2642927;
            12'd533: coeff = 24'd2652312;
            12'd534: coeff = 24'd2661710;
            12'd535: coeff = 24'd2671122;
            12'd536: coeff = 24'd2680547;
            12'd537: coeff = 24'd2689985;
            12'd538: coeff = 24'd2699437;
            12'd539: coeff = 24'd2708903;
            12'd540: coeff = 24'd2718381;
            12'd541: coeff = 24'd2727873;
            12'd542: coeff = 24'd2737379;
            12'd543: coeff = 24'd2746897;
            12'd544: coeff = 24'd2756429;
            12'd545: coeff = 24'd2765975;
            12'd546: coeff = 24'd2775533;
            12'd547: coeff = 24'd2785105;
            12'd548: coeff = 24'd2794690;
            12'd549: coeff = 24'd2804288;
            12'd550: coeff = 24'd2813899;
            12'd551: coeff = 24'd2823523;
            12'd552: coeff = 24'd2833161;
            12'd553: coeff = 24'd2842811;
            12'd554: coeff = 24'd2852475;
            12'd555: coeff = 24'd2862151;
            12'd556: coeff = 24'd2871841;
            12'd557: coeff = 24'd2881544;
            12'd558: coeff = 24'd2891259;
            12'd559: coeff = 24'd2900988;
            12'd560: coeff = 24'd2910729;
            12'd561: coeff = 24'd2920483;
            12'd562: coeff = 24'd2930251;
            12'd563: coeff = 24'd2940031;
            12'd564: coeff = 24'd2949824;
            12'd565: coeff = 24'd2959629;
            12'd566: coeff = 24'd2969448;
            12'd567: coeff = 24'd2979279;
            12'd568: coeff = 24'd2989123;
            12'd569: coeff = 24'd2998980;
            12'd570: coeff = 24'd3008849;
            12'd571: coeff = 24'd3018731;
            12'd572: coeff = 24'd3028626;
            12'd573: coeff = 24'd3038533;
            12'd574: coeff = 24'd3048453;
            12'd575: coeff = 24'd3058385;
            12'd576: coeff = 24'd3068330;
            12'd577: coeff = 24'd3078288;
            12'd578: coeff = 24'd3088258;
            12'd579: coeff = 24'd3098240;
            12'd580: coeff = 24'd3108235;
            12'd581: coeff = 24'd3118243;
            12'd582: coeff = 24'd3128262;
            12'd583: coeff = 24'd3138295;
            12'd584: coeff = 24'd3148339;
            12'd585: coeff = 24'd3158396;
            12'd586: coeff = 24'd3168465;
            12'd587: coeff = 24'd3178547;
            12'd588: coeff = 24'd3188640;
            12'd589: coeff = 24'd3198746;
            12'd590: coeff = 24'd3208865;
            12'd591: coeff = 24'd3218995;
            12'd592: coeff = 24'd3229138;
            12'd593: coeff = 24'd3239292;
            12'd594: coeff = 24'd3249459;
            12'd595: coeff = 24'd3259638;
            12'd596: coeff = 24'd3269829;
            12'd597: coeff = 24'd3280032;
            12'd598: coeff = 24'd3290247;
            12'd599: coeff = 24'd3300474;
            12'd600: coeff = 24'd3310713;
            12'd601: coeff = 24'd3320964;
            12'd602: coeff = 24'd3331227;
            12'd603: coeff = 24'd3341502;
            12'd604: coeff = 24'd3351789;
            12'd605: coeff = 24'd3362088;
            12'd606: coeff = 24'd3372398;
            12'd607: coeff = 24'd3382720;
            12'd608: coeff = 24'd3393054;
            12'd609: coeff = 24'd3403400;
            12'd610: coeff = 24'd3413758;
            12'd611: coeff = 24'd3424127;
            12'd612: coeff = 24'd3434508;
            12'd613: coeff = 24'd3444900;
            12'd614: coeff = 24'd3455305;
            12'd615: coeff = 24'd3465720;
            12'd616: coeff = 24'd3476148;
            12'd617: coeff = 24'd3486587;
            12'd618: coeff = 24'd3497037;
            12'd619: coeff = 24'd3507499;
            12'd620: coeff = 24'd3517973;
            12'd621: coeff = 24'd3528458;
            12'd622: coeff = 24'd3538954;
            12'd623: coeff = 24'd3549462;
            12'd624: coeff = 24'd3559982;
            12'd625: coeff = 24'd3570512;
            12'd626: coeff = 24'd3581054;
            12'd627: coeff = 24'd3591607;
            12'd628: coeff = 24'd3602172;
            12'd629: coeff = 24'd3612748;
            12'd630: coeff = 24'd3623335;
            12'd631: coeff = 24'd3633933;
            12'd632: coeff = 24'd3644543;
            12'd633: coeff = 24'd3655164;
            12'd634: coeff = 24'd3665795;
            12'd635: coeff = 24'd3676438;
            12'd636: coeff = 24'd3687092;
            12'd637: coeff = 24'd3697757;
            12'd638: coeff = 24'd3708434;
            12'd639: coeff = 24'd3719121;
            12'd640: coeff = 24'd3729819;
            12'd641: coeff = 24'd3740528;
            12'd642: coeff = 24'd3751248;
            12'd643: coeff = 24'd3761979;
            12'd644: coeff = 24'd3772721;
            12'd645: coeff = 24'd3783474;
            12'd646: coeff = 24'd3794237;
            12'd647: coeff = 24'd3805012;
            12'd648: coeff = 24'd3815797;
            12'd649: coeff = 24'd3826593;
            12'd650: coeff = 24'd3837400;
            12'd651: coeff = 24'd3848217;
            12'd652: coeff = 24'd3859045;
            12'd653: coeff = 24'd3869884;
            12'd654: coeff = 24'd3880733;
            12'd655: coeff = 24'd3891593;
            12'd656: coeff = 24'd3902464;
            12'd657: coeff = 24'd3913345;
            12'd658: coeff = 24'd3924237;
            12'd659: coeff = 24'd3935139;
            12'd660: coeff = 24'd3946052;
            12'd661: coeff = 24'd3956975;
            12'd662: coeff = 24'd3967908;
            12'd663: coeff = 24'd3978852;
            12'd664: coeff = 24'd3989807;
            12'd665: coeff = 24'd4000772;
            12'd666: coeff = 24'd4011747;
            12'd667: coeff = 24'd4022732;
            12'd668: coeff = 24'd4033728;
            12'd669: coeff = 24'd4044734;
            12'd670: coeff = 24'd4055750;
            12'd671: coeff = 24'd4066776;
            12'd672: coeff = 24'd4077812;
            12'd673: coeff = 24'd4088859;
            12'd674: coeff = 24'd4099916;
            12'd675: coeff = 24'd4110983;
            12'd676: coeff = 24'd4122060;
            12'd677: coeff = 24'd4133147;
            12'd678: coeff = 24'd4144244;
            12'd679: coeff = 24'd4155351;
            12'd680: coeff = 24'd4166468;
            12'd681: coeff = 24'd4177595;
            12'd682: coeff = 24'd4188731;
            12'd683: coeff = 24'd4199878;
            12'd684: coeff = 24'd4211035;
            12'd685: coeff = 24'd4222201;
            12'd686: coeff = 24'd4233377;
            12'd687: coeff = 24'd4244563;
            12'd688: coeff = 24'd4255759;
            12'd689: coeff = 24'd4266964;
            12'd690: coeff = 24'd4278180;
            12'd691: coeff = 24'd4289405;
            12'd692: coeff = 24'd4300639;
            12'd693: coeff = 24'd4311883;
            12'd694: coeff = 24'd4323137;
            12'd695: coeff = 24'd4334400;
            12'd696: coeff = 24'd4345673;
            12'd697: coeff = 24'd4356955;
            12'd698: coeff = 24'd4368247;
            12'd699: coeff = 24'd4379549;
            12'd700: coeff = 24'd4390859;
            12'd701: coeff = 24'd4402179;
            12'd702: coeff = 24'd4413509;
            12'd703: coeff = 24'd4424848;
            12'd704: coeff = 24'd4436196;
            12'd705: coeff = 24'd4447554;
            12'd706: coeff = 24'd4458921;
            12'd707: coeff = 24'd4470297;
            12'd708: coeff = 24'd4481682;
            12'd709: coeff = 24'd4493076;
            12'd710: coeff = 24'd4504480;
            12'd711: coeff = 24'd4515893;
            12'd712: coeff = 24'd4527315;
            12'd713: coeff = 24'd4538746;
            12'd714: coeff = 24'd4550186;
            12'd715: coeff = 24'd4561635;
            12'd716: coeff = 24'd4573093;
            12'd717: coeff = 24'd4584560;
            12'd718: coeff = 24'd4596036;
            12'd719: coeff = 24'd4607521;
            12'd720: coeff = 24'd4619015;
            12'd721: coeff = 24'd4630518;
            12'd722: coeff = 24'd4642030;
            12'd723: coeff = 24'd4653550;
            12'd724: coeff = 24'd4665079;
            12'd725: coeff = 24'd4676617;
            12'd726: coeff = 24'd4688164;
            12'd727: coeff = 24'd4699720;
            12'd728: coeff = 24'd4711284;
            12'd729: coeff = 24'd4722857;
            12'd730: coeff = 24'd4734438;
            12'd731: coeff = 24'd4746028;
            12'd732: coeff = 24'd4757627;
            12'd733: coeff = 24'd4769234;
            12'd734: coeff = 24'd4780849;
            12'd735: coeff = 24'd4792474;
            12'd736: coeff = 24'd4804106;
            12'd737: coeff = 24'd4815747;
            12'd738: coeff = 24'd4827397;
            12'd739: coeff = 24'd4839055;
            12'd740: coeff = 24'd4850721;
            12'd741: coeff = 24'd4862395;
            12'd742: coeff = 24'd4874078;
            12'd743: coeff = 24'd4885769;
            12'd744: coeff = 24'd4897469;
            12'd745: coeff = 24'd4909176;
            12'd746: coeff = 24'd4920892;
            12'd747: coeff = 24'd4932616;
            12'd748: coeff = 24'd4944348;
            12'd749: coeff = 24'd4956088;
            12'd750: coeff = 24'd4967837;
            12'd751: coeff = 24'd4979593;
            12'd752: coeff = 24'd4991357;
            12'd753: coeff = 24'd5003130;
            12'd754: coeff = 24'd5014910;
            12'd755: coeff = 24'd5026698;
            12'd756: coeff = 24'd5038495;
            12'd757: coeff = 24'd5050299;
            12'd758: coeff = 24'd5062111;
            12'd759: coeff = 24'd5073930;
            12'd760: coeff = 24'd5085758;
            12'd761: coeff = 24'd5097593;
            12'd762: coeff = 24'd5109436;
            12'd763: coeff = 24'd5121287;
            12'd764: coeff = 24'd5133146;
            12'd765: coeff = 24'd5145012;
            12'd766: coeff = 24'd5156886;
            12'd767: coeff = 24'd5168767;
            12'd768: coeff = 24'd5180656;
            12'd769: coeff = 24'd5192552;
            12'd770: coeff = 24'd5204457;
            12'd771: coeff = 24'd5216368;
            12'd772: coeff = 24'd5228287;
            12'd773: coeff = 24'd5240214;
            12'd774: coeff = 24'd5252147;
            12'd775: coeff = 24'd5264089;
            12'd776: coeff = 24'd5276037;
            12'd777: coeff = 24'd5287993;
            12'd778: coeff = 24'd5299957;
            12'd779: coeff = 24'd5311927;
            12'd780: coeff = 24'd5323905;
            12'd781: coeff = 24'd5335890;
            12'd782: coeff = 24'd5347882;
            12'd783: coeff = 24'd5359881;
            12'd784: coeff = 24'd5371888;
            12'd785: coeff = 24'd5383901;
            12'd786: coeff = 24'd5395922;
            12'd787: coeff = 24'd5407950;
            12'd788: coeff = 24'd5419984;
            12'd789: coeff = 24'd5432026;
            12'd790: coeff = 24'd5444075;
            12'd791: coeff = 24'd5456130;
            12'd792: coeff = 24'd5468193;
            12'd793: coeff = 24'd5480262;
            12'd794: coeff = 24'd5492338;
            12'd795: coeff = 24'd5504421;
            12'd796: coeff = 24'd5516511;
            12'd797: coeff = 24'd5528608;
            12'd798: coeff = 24'd5540711;
            12'd799: coeff = 24'd5552821;
            12'd800: coeff = 24'd5564938;
            12'd801: coeff = 24'd5577061;
            12'd802: coeff = 24'd5589191;
            12'd803: coeff = 24'd5601327;
            12'd804: coeff = 24'd5613471;
            12'd805: coeff = 24'd5625620;
            12'd806: coeff = 24'd5637776;
            12'd807: coeff = 24'd5649939;
            12'd808: coeff = 24'd5662108;
            12'd809: coeff = 24'd5674284;
            12'd810: coeff = 24'd5686465;
            12'd811: coeff = 24'd5698654;
            12'd812: coeff = 24'd5710848;
            12'd813: coeff = 24'd5723049;
            12'd814: coeff = 24'd5735256;
            12'd815: coeff = 24'd5747470;
            12'd816: coeff = 24'd5759689;
            12'd817: coeff = 24'd5771915;
            12'd818: coeff = 24'd5784147;
            12'd819: coeff = 24'd5796385;
            12'd820: coeff = 24'd5808629;
            12'd821: coeff = 24'd5820880;
            12'd822: coeff = 24'd5833136;
            12'd823: coeff = 24'd5845398;
            12'd824: coeff = 24'd5857666;
            12'd825: coeff = 24'd5869941;
            12'd826: coeff = 24'd5882221;
            12'd827: coeff = 24'd5894507;
            12'd828: coeff = 24'd5906799;
            12'd829: coeff = 24'd5919097;
            12'd830: coeff = 24'd5931401;
            12'd831: coeff = 24'd5943710;
            12'd832: coeff = 24'd5956025;
            12'd833: coeff = 24'd5968346;
            12'd834: coeff = 24'd5980673;
            12'd835: coeff = 24'd5993005;
            12'd836: coeff = 24'd6005343;
            12'd837: coeff = 24'd6017686;
            12'd838: coeff = 24'd6030035;
            12'd839: coeff = 24'd6042390;
            12'd840: coeff = 24'd6054750;
            12'd841: coeff = 24'd6067116;
            12'd842: coeff = 24'd6079487;
            12'd843: coeff = 24'd6091864;
            12'd844: coeff = 24'd6104246;
            12'd845: coeff = 24'd6116633;
            12'd846: coeff = 24'd6129026;
            12'd847: coeff = 24'd6141424;
            12'd848: coeff = 24'd6153827;
            12'd849: coeff = 24'd6166236;
            12'd850: coeff = 24'd6178649;
            12'd851: coeff = 24'd6191068;
            12'd852: coeff = 24'd6203493;
            12'd853: coeff = 24'd6215922;
            12'd854: coeff = 24'd6228356;
            12'd855: coeff = 24'd6240796;
            12'd856: coeff = 24'd6253241;
            12'd857: coeff = 24'd6265690;
            12'd858: coeff = 24'd6278145;
            12'd859: coeff = 24'd6290604;
            12'd860: coeff = 24'd6303069;
            12'd861: coeff = 24'd6315538;
            12'd862: coeff = 24'd6328013;
            12'd863: coeff = 24'd6340492;
            12'd864: coeff = 24'd6352976;
            12'd865: coeff = 24'd6365465;
            12'd866: coeff = 24'd6377958;
            12'd867: coeff = 24'd6390456;
            12'd868: coeff = 24'd6402959;
            12'd869: coeff = 24'd6415467;
            12'd870: coeff = 24'd6427979;
            12'd871: coeff = 24'd6440496;
            12'd872: coeff = 24'd6453018;
            12'd873: coeff = 24'd6465544;
            12'd874: coeff = 24'd6478074;
            12'd875: coeff = 24'd6490609;
            12'd876: coeff = 24'd6503149;
            12'd877: coeff = 24'd6515693;
            12'd878: coeff = 24'd6528241;
            12'd879: coeff = 24'd6540794;
            12'd880: coeff = 24'd6553351;
            12'd881: coeff = 24'd6565913;
            12'd882: coeff = 24'd6578478;
            12'd883: coeff = 24'd6591048;
            12'd884: coeff = 24'd6603623;
            12'd885: coeff = 24'd6616201;
            12'd886: coeff = 24'd6628784;
            12'd887: coeff = 24'd6641370;
            12'd888: coeff = 24'd6653961;
            12'd889: coeff = 24'd6666556;
            12'd890: coeff = 24'd6679155;
            12'd891: coeff = 24'd6691758;
            12'd892: coeff = 24'd6704365;
            12'd893: coeff = 24'd6716976;
            12'd894: coeff = 24'd6729591;
            12'd895: coeff = 24'd6742210;
            12'd896: coeff = 24'd6754833;
            12'd897: coeff = 24'd6767459;
            12'd898: coeff = 24'd6780090;
            12'd899: coeff = 24'd6792724;
            12'd900: coeff = 24'd6805362;
            12'd901: coeff = 24'd6818003;
            12'd902: coeff = 24'd6830649;
            12'd903: coeff = 24'd6843298;
            12'd904: coeff = 24'd6855950;
            12'd905: coeff = 24'd6868607;
            12'd906: coeff = 24'd6881267;
            12'd907: coeff = 24'd6893930;
            12'd908: coeff = 24'd6906597;
            12'd909: coeff = 24'd6919267;
            12'd910: coeff = 24'd6931941;
            12'd911: coeff = 24'd6944618;
            12'd912: coeff = 24'd6957299;
            12'd913: coeff = 24'd6969983;
            12'd914: coeff = 24'd6982670;
            12'd915: coeff = 24'd6995361;
            12'd916: coeff = 24'd7008055;
            12'd917: coeff = 24'd7020752;
            12'd918: coeff = 24'd7033453;
            12'd919: coeff = 24'd7046156;
            12'd920: coeff = 24'd7058863;
            12'd921: coeff = 24'd7071573;
            12'd922: coeff = 24'd7084286;
            12'd923: coeff = 24'd7097002;
            12'd924: coeff = 24'd7109721;
            12'd925: coeff = 24'd7122443;
            12'd926: coeff = 24'd7135169;
            12'd927: coeff = 24'd7147897;
            12'd928: coeff = 24'd7160628;
            12'd929: coeff = 24'd7173362;
            12'd930: coeff = 24'd7186098;
            12'd931: coeff = 24'd7198838;
            12'd932: coeff = 24'd7211580;
            12'd933: coeff = 24'd7224325;
            12'd934: coeff = 24'd7237073;
            12'd935: coeff = 24'd7249824;
            12'd936: coeff = 24'd7262577;
            12'd937: coeff = 24'd7275333;
            12'd938: coeff = 24'd7288092;
            12'd939: coeff = 24'd7300853;
            12'd940: coeff = 24'd7313617;
            12'd941: coeff = 24'd7326383;
            12'd942: coeff = 24'd7339152;
            12'd943: coeff = 24'd7351923;
            12'd944: coeff = 24'd7364696;
            12'd945: coeff = 24'd7377473;
            12'd946: coeff = 24'd7390251;
            12'd947: coeff = 24'd7403032;
            12'd948: coeff = 24'd7415815;
            12'd949: coeff = 24'd7428600;
            12'd950: coeff = 24'd7441388;
            12'd951: coeff = 24'd7454178;
            12'd952: coeff = 24'd7466970;
            12'd953: coeff = 24'd7479764;
            12'd954: coeff = 24'd7492561;
            12'd955: coeff = 24'd7505359;
            12'd956: coeff = 24'd7518160;
            12'd957: coeff = 24'd7530962;
            12'd958: coeff = 24'd7543767;
            12'd959: coeff = 24'd7556574;
            12'd960: coeff = 24'd7569382;
            12'd961: coeff = 24'd7582193;
            12'd962: coeff = 24'd7595005;
            12'd963: coeff = 24'd7607820;
            12'd964: coeff = 24'd7620636;
            12'd965: coeff = 24'd7633454;
            12'd966: coeff = 24'd7646273;
            12'd967: coeff = 24'd7659095;
            12'd968: coeff = 24'd7671918;
            12'd969: coeff = 24'd7684743;
            12'd970: coeff = 24'd7697570;
            12'd971: coeff = 24'd7710398;
            12'd972: coeff = 24'd7723227;
            12'd973: coeff = 24'd7736059;
            12'd974: coeff = 24'd7748892;
            12'd975: coeff = 24'd7761726;
            12'd976: coeff = 24'd7774562;
            12'd977: coeff = 24'd7787399;
            12'd978: coeff = 24'd7800238;
            12'd979: coeff = 24'd7813078;
            12'd980: coeff = 24'd7825919;
            12'd981: coeff = 24'd7838762;
            12'd982: coeff = 24'd7851606;
            12'd983: coeff = 24'd7864452;
            12'd984: coeff = 24'd7877298;
            12'd985: coeff = 24'd7890146;
            12'd986: coeff = 24'd7902995;
            12'd987: coeff = 24'd7915845;
            12'd988: coeff = 24'd7928696;
            12'd989: coeff = 24'd7941548;
            12'd990: coeff = 24'd7954402;
            12'd991: coeff = 24'd7967256;
            12'd992: coeff = 24'd7980112;
            12'd993: coeff = 24'd7992968;
            12'd994: coeff = 24'd8005825;
            12'd995: coeff = 24'd8018683;
            12'd996: coeff = 24'd8031542;
            12'd997: coeff = 24'd8044402;
            12'd998: coeff = 24'd8057263;
            12'd999: coeff = 24'd8070124;
            12'd1000: coeff = 24'd8082986;
            12'd1001: coeff = 24'd8095849;
            12'd1002: coeff = 24'd8108713;
            12'd1003: coeff = 24'd8121577;
            12'd1004: coeff = 24'd8134442;
            12'd1005: coeff = 24'd8147308;
            12'd1006: coeff = 24'd8160174;
            12'd1007: coeff = 24'd8173040;
            12'd1008: coeff = 24'd8185907;
            12'd1009: coeff = 24'd8198775;
            12'd1010: coeff = 24'd8211643;
            12'd1011: coeff = 24'd8224511;
            12'd1012: coeff = 24'd8237380;
            12'd1013: coeff = 24'd8250249;
            12'd1014: coeff = 24'd8263119;
            12'd1015: coeff = 24'd8275989;
            12'd1016: coeff = 24'd8288859;
            12'd1017: coeff = 24'd8301729;
            12'd1018: coeff = 24'd8314600;
            12'd1019: coeff = 24'd8327470;
            12'd1020: coeff = 24'd8340341;
            12'd1021: coeff = 24'd8353212;
            12'd1022: coeff = 24'd8366083;
            12'd1023: coeff = 24'd8378954;
            12'd1024: coeff = 24'd8391825;
            12'd1025: coeff = 24'd8404696;
            12'd1026: coeff = 24'd8417567;
            12'd1027: coeff = 24'd8430438;
            12'd1028: coeff = 24'd8443309;
            12'd1029: coeff = 24'd8456180;
            12'd1030: coeff = 24'd8469051;
            12'd1031: coeff = 24'd8481921;
            12'd1032: coeff = 24'd8494791;
            12'd1033: coeff = 24'd8507661;
            12'd1034: coeff = 24'd8520531;
            12'd1035: coeff = 24'd8533400;
            12'd1036: coeff = 24'd8546269;
            12'd1037: coeff = 24'd8559138;
            12'd1038: coeff = 24'd8572006;
            12'd1039: coeff = 24'd8584874;
            12'd1040: coeff = 24'd8597741;
            12'd1041: coeff = 24'd8610608;
            12'd1042: coeff = 24'd8623474;
            12'd1043: coeff = 24'd8636340;
            12'd1044: coeff = 24'd8649205;
            12'd1045: coeff = 24'd8662070;
            12'd1046: coeff = 24'd8674934;
            12'd1047: coeff = 24'd8687797;
            12'd1048: coeff = 24'd8700660;
            12'd1049: coeff = 24'd8713522;
            12'd1050: coeff = 24'd8726383;
            12'd1051: coeff = 24'd8739243;
            12'd1052: coeff = 24'd8752102;
            12'd1053: coeff = 24'd8764961;
            12'd1054: coeff = 24'd8777819;
            12'd1055: coeff = 24'd8790675;
            12'd1056: coeff = 24'd8803531;
            12'd1057: coeff = 24'd8816386;
            12'd1058: coeff = 24'd8829240;
            12'd1059: coeff = 24'd8842093;
            12'd1060: coeff = 24'd8854945;
            12'd1061: coeff = 24'd8867795;
            12'd1062: coeff = 24'd8880645;
            12'd1063: coeff = 24'd8893493;
            12'd1064: coeff = 24'd8906340;
            12'd1065: coeff = 24'd8919186;
            12'd1066: coeff = 24'd8932031;
            12'd1067: coeff = 24'd8944874;
            12'd1068: coeff = 24'd8957716;
            12'd1069: coeff = 24'd8970557;
            12'd1070: coeff = 24'd8983397;
            12'd1071: coeff = 24'd8996235;
            12'd1072: coeff = 24'd9009071;
            12'd1073: coeff = 24'd9021906;
            12'd1074: coeff = 24'd9034740;
            12'd1075: coeff = 24'd9047572;
            12'd1076: coeff = 24'd9060403;
            12'd1077: coeff = 24'd9073232;
            12'd1078: coeff = 24'd9086059;
            12'd1079: coeff = 24'd9098885;
            12'd1080: coeff = 24'd9111709;
            12'd1081: coeff = 24'd9124531;
            12'd1082: coeff = 24'd9137352;
            12'd1083: coeff = 24'd9150170;
            12'd1084: coeff = 24'd9162988;
            12'd1085: coeff = 24'd9175803;
            12'd1086: coeff = 24'd9188616;
            12'd1087: coeff = 24'd9201428;
            12'd1088: coeff = 24'd9214237;
            12'd1089: coeff = 24'd9227045;
            12'd1090: coeff = 24'd9239851;
            12'd1091: coeff = 24'd9252654;
            12'd1092: coeff = 24'd9265456;
            12'd1093: coeff = 24'd9278255;
            12'd1094: coeff = 24'd9291053;
            12'd1095: coeff = 24'd9303848;
            12'd1096: coeff = 24'd9316641;
            12'd1097: coeff = 24'd9329432;
            12'd1098: coeff = 24'd9342221;
            12'd1099: coeff = 24'd9355008;
            12'd1100: coeff = 24'd9367792;
            12'd1101: coeff = 24'd9380574;
            12'd1102: coeff = 24'd9393354;
            12'd1103: coeff = 24'd9406131;
            12'd1104: coeff = 24'd9418906;
            12'd1105: coeff = 24'd9431678;
            12'd1106: coeff = 24'd9444448;
            12'd1107: coeff = 24'd9457216;
            12'd1108: coeff = 24'd9469981;
            12'd1109: coeff = 24'd9482743;
            12'd1110: coeff = 24'd9495503;
            12'd1111: coeff = 24'd9508260;
            12'd1112: coeff = 24'd9521015;
            12'd1113: coeff = 24'd9533767;
            12'd1114: coeff = 24'd9546516;
            12'd1115: coeff = 24'd9559262;
            12'd1116: coeff = 24'd9572006;
            12'd1117: coeff = 24'd9584747;
            12'd1118: coeff = 24'd9597485;
            12'd1119: coeff = 24'd9610221;
            12'd1120: coeff = 24'd9622953;
            12'd1121: coeff = 24'd9635683;
            12'd1122: coeff = 24'd9648409;
            12'd1123: coeff = 24'd9661133;
            12'd1124: coeff = 24'd9673854;
            12'd1125: coeff = 24'd9686571;
            12'd1126: coeff = 24'd9699286;
            12'd1127: coeff = 24'd9711997;
            12'd1128: coeff = 24'd9724706;
            12'd1129: coeff = 24'd9737411;
            12'd1130: coeff = 24'd9750113;
            12'd1131: coeff = 24'd9762812;
            12'd1132: coeff = 24'd9775507;
            12'd1133: coeff = 24'd9788200;
            12'd1134: coeff = 24'd9800889;
            12'd1135: coeff = 24'd9813574;
            12'd1136: coeff = 24'd9826257;
            12'd1137: coeff = 24'd9838936;
            12'd1138: coeff = 24'd9851611;
            12'd1139: coeff = 24'd9864283;
            12'd1140: coeff = 24'd9876952;
            12'd1141: coeff = 24'd9889617;
            12'd1142: coeff = 24'd9902279;
            12'd1143: coeff = 24'd9914937;
            12'd1144: coeff = 24'd9927591;
            12'd1145: coeff = 24'd9940242;
            12'd1146: coeff = 24'd9952889;
            12'd1147: coeff = 24'd9965533;
            12'd1148: coeff = 24'd9978173;
            12'd1149: coeff = 24'd9990809;
            12'd1150: coeff = 24'd10003441;
            12'd1151: coeff = 24'd10016069;
            12'd1152: coeff = 24'd10028694;
            12'd1153: coeff = 24'd10041315;
            12'd1154: coeff = 24'd10053932;
            12'd1155: coeff = 24'd10066545;
            12'd1156: coeff = 24'd10079154;
            12'd1157: coeff = 24'd10091759;
            12'd1158: coeff = 24'd10104360;
            12'd1159: coeff = 24'd10116957;
            12'd1160: coeff = 24'd10129550;
            12'd1161: coeff = 24'd10142138;
            12'd1162: coeff = 24'd10154723;
            12'd1163: coeff = 24'd10167304;
            12'd1164: coeff = 24'd10179880;
            12'd1165: coeff = 24'd10192452;
            12'd1166: coeff = 24'd10205020;
            12'd1167: coeff = 24'd10217584;
            12'd1168: coeff = 24'd10230143;
            12'd1169: coeff = 24'd10242698;
            12'd1170: coeff = 24'd10255248;
            12'd1171: coeff = 24'd10267795;
            12'd1172: coeff = 24'd10280336;
            12'd1173: coeff = 24'd10292874;
            12'd1174: coeff = 24'd10305407;
            12'd1175: coeff = 24'd10317935;
            12'd1176: coeff = 24'd10330459;
            12'd1177: coeff = 24'd10342978;
            12'd1178: coeff = 24'd10355492;
            12'd1179: coeff = 24'd10368002;
            12'd1180: coeff = 24'd10380508;
            12'd1181: coeff = 24'd10393008;
            12'd1182: coeff = 24'd10405504;
            12'd1183: coeff = 24'd10417995;
            12'd1184: coeff = 24'd10430482;
            12'd1185: coeff = 24'd10442963;
            12'd1186: coeff = 24'd10455440;
            12'd1187: coeff = 24'd10467912;
            12'd1188: coeff = 24'd10480379;
            12'd1189: coeff = 24'd10492841;
            12'd1190: coeff = 24'd10505298;
            12'd1191: coeff = 24'd10517750;
            12'd1192: coeff = 24'd10530197;
            12'd1193: coeff = 24'd10542639;
            12'd1194: coeff = 24'd10555076;
            12'd1195: coeff = 24'd10567508;
            12'd1196: coeff = 24'd10579935;
            12'd1197: coeff = 24'd10592357;
            12'd1198: coeff = 24'd10604773;
            12'd1199: coeff = 24'd10617184;
            12'd1200: coeff = 24'd10629590;
            12'd1201: coeff = 24'd10641991;
            12'd1202: coeff = 24'd10654386;
            12'd1203: coeff = 24'd10666776;
            12'd1204: coeff = 24'd10679161;
            12'd1205: coeff = 24'd10691540;
            12'd1206: coeff = 24'd10703914;
            12'd1207: coeff = 24'd10716283;
            12'd1208: coeff = 24'd10728646;
            12'd1209: coeff = 24'd10741003;
            12'd1210: coeff = 24'd10753355;
            12'd1211: coeff = 24'd10765701;
            12'd1212: coeff = 24'd10778042;
            12'd1213: coeff = 24'd10790377;
            12'd1214: coeff = 24'd10802706;
            12'd1215: coeff = 24'd10815030;
            12'd1216: coeff = 24'd10827348;
            12'd1217: coeff = 24'd10839660;
            12'd1218: coeff = 24'd10851967;
            12'd1219: coeff = 24'd10864268;
            12'd1220: coeff = 24'd10876563;
            12'd1221: coeff = 24'd10888852;
            12'd1222: coeff = 24'd10901135;
            12'd1223: coeff = 24'd10913412;
            12'd1224: coeff = 24'd10925683;
            12'd1225: coeff = 24'd10937949;
            12'd1226: coeff = 24'd10950208;
            12'd1227: coeff = 24'd10962461;
            12'd1228: coeff = 24'd10974709;
            12'd1229: coeff = 24'd10986950;
            12'd1230: coeff = 24'd10999185;
            12'd1231: coeff = 24'd11011414;
            12'd1232: coeff = 24'd11023636;
            12'd1233: coeff = 24'd11035853;
            12'd1234: coeff = 24'd11048063;
            12'd1235: coeff = 24'd11060267;
            12'd1236: coeff = 24'd11072465;
            12'd1237: coeff = 24'd11084656;
            12'd1238: coeff = 24'd11096841;
            12'd1239: coeff = 24'd11109020;
            12'd1240: coeff = 24'd11121192;
            12'd1241: coeff = 24'd11133358;
            12'd1242: coeff = 24'd11145518;
            12'd1243: coeff = 24'd11157670;
            12'd1244: coeff = 24'd11169817;
            12'd1245: coeff = 24'd11181957;
            12'd1246: coeff = 24'd11194090;
            12'd1247: coeff = 24'd11206217;
            12'd1248: coeff = 24'd11218337;
            12'd1249: coeff = 24'd11230450;
            12'd1250: coeff = 24'd11242557;
            12'd1251: coeff = 24'd11254656;
            12'd1252: coeff = 24'd11266750;
            12'd1253: coeff = 24'd11278836;
            12'd1254: coeff = 24'd11290916;
            12'd1255: coeff = 24'd11302988;
            12'd1256: coeff = 24'd11315054;
            12'd1257: coeff = 24'd11327113;
            12'd1258: coeff = 24'd11339166;
            12'd1259: coeff = 24'd11351211;
            12'd1260: coeff = 24'd11363249;
            12'd1261: coeff = 24'd11375280;
            12'd1262: coeff = 24'd11387304;
            12'd1263: coeff = 24'd11399321;
            12'd1264: coeff = 24'd11411331;
            12'd1265: coeff = 24'd11423334;
            12'd1266: coeff = 24'd11435330;
            12'd1267: coeff = 24'd11447319;
            12'd1268: coeff = 24'd11459300;
            12'd1269: coeff = 24'd11471274;
            12'd1270: coeff = 24'd11483241;
            12'd1271: coeff = 24'd11495201;
            12'd1272: coeff = 24'd11507153;
            12'd1273: coeff = 24'd11519098;
            12'd1274: coeff = 24'd11531035;
            12'd1275: coeff = 24'd11542966;
            12'd1276: coeff = 24'd11554888;
            12'd1277: coeff = 24'd11566804;
            12'd1278: coeff = 24'd11578711;
            12'd1279: coeff = 24'd11590612;
            12'd1280: coeff = 24'd11602504;
            12'd1281: coeff = 24'd11614390;
            12'd1282: coeff = 24'd11626267;
            12'd1283: coeff = 24'd11638137;
            12'd1284: coeff = 24'd11650000;
            12'd1285: coeff = 24'd11661854;
            12'd1286: coeff = 24'd11673701;
            12'd1287: coeff = 24'd11685540;
            12'd1288: coeff = 24'd11697372;
            12'd1289: coeff = 24'd11709196;
            12'd1290: coeff = 24'd11721011;
            12'd1291: coeff = 24'd11732819;
            12'd1292: coeff = 24'd11744620;
            12'd1293: coeff = 24'd11756412;
            12'd1294: coeff = 24'd11768196;
            12'd1295: coeff = 24'd11779972;
            12'd1296: coeff = 24'd11791741;
            12'd1297: coeff = 24'd11803501;
            12'd1298: coeff = 24'd11815253;
            12'd1299: coeff = 24'd11826998;
            12'd1300: coeff = 24'd11838734;
            12'd1301: coeff = 24'd11850462;
            12'd1302: coeff = 24'd11862182;
            12'd1303: coeff = 24'd11873893;
            12'd1304: coeff = 24'd11885597;
            12'd1305: coeff = 24'd11897292;
            12'd1306: coeff = 24'd11908979;
            12'd1307: coeff = 24'd11920658;
            12'd1308: coeff = 24'd11932328;
            12'd1309: coeff = 24'd11943990;
            12'd1310: coeff = 24'd11955644;
            12'd1311: coeff = 24'd11967289;
            12'd1312: coeff = 24'd11978926;
            12'd1313: coeff = 24'd11990554;
            12'd1314: coeff = 24'd12002174;
            12'd1315: coeff = 24'd12013786;
            12'd1316: coeff = 24'd12025389;
            12'd1317: coeff = 24'd12036983;
            12'd1318: coeff = 24'd12048569;
            12'd1319: coeff = 24'd12060146;
            12'd1320: coeff = 24'd12071714;
            12'd1321: coeff = 24'd12083274;
            12'd1322: coeff = 24'd12094825;
            12'd1323: coeff = 24'd12106368;
            12'd1324: coeff = 24'd12117901;
            12'd1325: coeff = 24'd12129426;
            12'd1326: coeff = 24'd12140942;
            12'd1327: coeff = 24'd12152449;
            12'd1328: coeff = 24'd12163948;
            12'd1329: coeff = 24'd12175437;
            12'd1330: coeff = 24'd12186918;
            12'd1331: coeff = 24'd12198389;
            12'd1332: coeff = 24'd12209852;
            12'd1333: coeff = 24'd12221306;
            12'd1334: coeff = 24'd12232750;
            12'd1335: coeff = 24'd12244186;
            12'd1336: coeff = 24'd12255612;
            12'd1337: coeff = 24'd12267030;
            12'd1338: coeff = 24'd12278438;
            12'd1339: coeff = 24'd12289837;
            12'd1340: coeff = 24'd12301227;
            12'd1341: coeff = 24'd12312608;
            12'd1342: coeff = 24'd12323979;
            12'd1343: coeff = 24'd12335341;
            12'd1344: coeff = 24'd12346694;
            12'd1345: coeff = 24'd12358038;
            12'd1346: coeff = 24'd12369372;
            12'd1347: coeff = 24'd12380697;
            12'd1348: coeff = 24'd12392012;
            12'd1349: coeff = 24'd12403318;
            12'd1350: coeff = 24'd12414615;
            12'd1351: coeff = 24'd12425902;
            12'd1352: coeff = 24'd12437180;
            12'd1353: coeff = 24'd12448448;
            12'd1354: coeff = 24'd12459706;
            12'd1355: coeff = 24'd12470955;
            12'd1356: coeff = 24'd12482194;
            12'd1357: coeff = 24'd12493424;
            12'd1358: coeff = 24'd12504644;
            12'd1359: coeff = 24'd12515854;
            12'd1360: coeff = 24'd12527055;
            12'd1361: coeff = 24'd12538246;
            12'd1362: coeff = 24'd12549427;
            12'd1363: coeff = 24'd12560598;
            12'd1364: coeff = 24'd12571760;
            12'd1365: coeff = 24'd12582911;
            12'd1366: coeff = 24'd12594053;
            12'd1367: coeff = 24'd12605185;
            12'd1368: coeff = 24'd12616307;
            12'd1369: coeff = 24'd12627419;
            12'd1370: coeff = 24'd12638521;
            12'd1371: coeff = 24'd12649613;
            12'd1372: coeff = 24'd12660695;
            12'd1373: coeff = 24'd12671767;
            12'd1374: coeff = 24'd12682829;
            12'd1375: coeff = 24'd12693880;
            12'd1376: coeff = 24'd12704922;
            12'd1377: coeff = 24'd12715953;
            12'd1378: coeff = 24'd12726975;
            12'd1379: coeff = 24'd12737986;
            12'd1380: coeff = 24'd12748986;
            12'd1381: coeff = 24'd12759977;
            12'd1382: coeff = 24'd12770957;
            12'd1383: coeff = 24'd12781927;
            12'd1384: coeff = 24'd12792887;
            12'd1385: coeff = 24'd12803836;
            12'd1386: coeff = 24'd12814775;
            12'd1387: coeff = 24'd12825703;
            12'd1388: coeff = 24'd12836621;
            12'd1389: coeff = 24'd12847528;
            12'd1390: coeff = 24'd12858425;
            12'd1391: coeff = 24'd12869312;
            12'd1392: coeff = 24'd12880188;
            12'd1393: coeff = 24'd12891053;
            12'd1394: coeff = 24'd12901908;
            12'd1395: coeff = 24'd12912752;
            12'd1396: coeff = 24'd12923585;
            12'd1397: coeff = 24'd12934408;
            12'd1398: coeff = 24'd12945220;
            12'd1399: coeff = 24'd12956021;
            12'd1400: coeff = 24'd12966812;
            12'd1401: coeff = 24'd12977592;
            12'd1402: coeff = 24'd12988361;
            12'd1403: coeff = 24'd12999119;
            12'd1404: coeff = 24'd13009866;
            12'd1405: coeff = 24'd13020603;
            12'd1406: coeff = 24'd13031328;
            12'd1407: coeff = 24'd13042043;
            12'd1408: coeff = 24'd13052747;
            12'd1409: coeff = 24'd13063439;
            12'd1410: coeff = 24'd13074121;
            12'd1411: coeff = 24'd13084791;
            12'd1412: coeff = 24'd13095451;
            12'd1413: coeff = 24'd13106100;
            12'd1414: coeff = 24'd13116737;
            12'd1415: coeff = 24'd13127363;
            12'd1416: coeff = 24'd13137978;
            12'd1417: coeff = 24'd13148582;
            12'd1418: coeff = 24'd13159175;
            12'd1419: coeff = 24'd13169756;
            12'd1420: coeff = 24'd13180327;
            12'd1421: coeff = 24'd13190886;
            12'd1422: coeff = 24'd13201433;
            12'd1423: coeff = 24'd13211970;
            12'd1424: coeff = 24'd13222494;
            12'd1425: coeff = 24'd13233008;
            12'd1426: coeff = 24'd13243510;
            12'd1427: coeff = 24'd13254001;
            12'd1428: coeff = 24'd13264480;
            12'd1429: coeff = 24'd13274948;
            12'd1430: coeff = 24'd13285404;
            12'd1431: coeff = 24'd13295849;
            12'd1432: coeff = 24'd13306282;
            12'd1433: coeff = 24'd13316704;
            12'd1434: coeff = 24'd13327114;
            12'd1435: coeff = 24'd13337512;
            12'd1436: coeff = 24'd13347899;
            12'd1437: coeff = 24'd13358274;
            12'd1438: coeff = 24'd13368638;
            12'd1439: coeff = 24'd13378989;
            12'd1440: coeff = 24'd13389329;
            12'd1441: coeff = 24'd13399657;
            12'd1442: coeff = 24'd13409974;
            12'd1443: coeff = 24'd13420278;
            12'd1444: coeff = 24'd13430571;
            12'd1445: coeff = 24'd13440852;
            12'd1446: coeff = 24'd13451121;
            12'd1447: coeff = 24'd13461378;
            12'd1448: coeff = 24'd13471623;
            12'd1449: coeff = 24'd13481856;
            12'd1450: coeff = 24'd13492077;
            12'd1451: coeff = 24'd13502286;
            12'd1452: coeff = 24'd13512483;
            12'd1453: coeff = 24'd13522668;
            12'd1454: coeff = 24'd13532841;
            12'd1455: coeff = 24'd13543002;
            12'd1456: coeff = 24'd13553150;
            12'd1457: coeff = 24'd13563287;
            12'd1458: coeff = 24'd13573411;
            12'd1459: coeff = 24'd13583523;
            12'd1460: coeff = 24'd13593623;
            12'd1461: coeff = 24'd13603711;
            12'd1462: coeff = 24'd13613786;
            12'd1463: coeff = 24'd13623849;
            12'd1464: coeff = 24'd13633900;
            12'd1465: coeff = 24'd13643938;
            12'd1466: coeff = 24'd13653964;
            12'd1467: coeff = 24'd13663978;
            12'd1468: coeff = 24'd13673979;
            12'd1469: coeff = 24'd13683968;
            12'd1470: coeff = 24'd13693944;
            12'd1471: coeff = 24'd13703908;
            12'd1472: coeff = 24'd13713859;
            12'd1473: coeff = 24'd13723798;
            12'd1474: coeff = 24'd13733724;
            12'd1475: coeff = 24'd13743637;
            12'd1476: coeff = 24'd13753538;
            12'd1477: coeff = 24'd13763427;
            12'd1478: coeff = 24'd13773302;
            12'd1479: coeff = 24'd13783165;
            12'd1480: coeff = 24'd13793016;
            12'd1481: coeff = 24'd13802853;
            12'd1482: coeff = 24'd13812678;
            12'd1483: coeff = 24'd13822490;
            12'd1484: coeff = 24'd13832289;
            12'd1485: coeff = 24'd13842076;
            12'd1486: coeff = 24'd13851850;
            12'd1487: coeff = 24'd13861610;
            12'd1488: coeff = 24'd13871358;
            12'd1489: coeff = 24'd13881093;
            12'd1490: coeff = 24'd13890815;
            12'd1491: coeff = 24'd13900524;
            12'd1492: coeff = 24'd13910220;
            12'd1493: coeff = 24'd13919903;
            12'd1494: coeff = 24'd13929574;
            12'd1495: coeff = 24'd13939231;
            12'd1496: coeff = 24'd13948875;
            12'd1497: coeff = 24'd13958505;
            12'd1498: coeff = 24'd13968123;
            12'd1499: coeff = 24'd13977728;
            12'd1500: coeff = 24'd13987319;
            12'd1501: coeff = 24'd13996898;
            12'd1502: coeff = 24'd14006463;
            12'd1503: coeff = 24'd14016015;
            12'd1504: coeff = 24'd14025553;
            12'd1505: coeff = 24'd14035079;
            12'd1506: coeff = 24'd14044591;
            12'd1507: coeff = 24'd14054089;
            12'd1508: coeff = 24'd14063575;
            12'd1509: coeff = 24'd14073047;
            12'd1510: coeff = 24'd14082505;
            12'd1511: coeff = 24'd14091951;
            12'd1512: coeff = 24'd14101383;
            12'd1513: coeff = 24'd14110801;
            12'd1514: coeff = 24'd14120206;
            12'd1515: coeff = 24'd14129597;
            12'd1516: coeff = 24'd14138975;
            12'd1517: coeff = 24'd14148340;
            12'd1518: coeff = 24'd14157690;
            12'd1519: coeff = 24'd14167028;
            12'd1520: coeff = 24'd14176351;
            12'd1521: coeff = 24'd14185661;
            12'd1522: coeff = 24'd14194958;
            12'd1523: coeff = 24'd14204240;
            12'd1524: coeff = 24'd14213509;
            12'd1525: coeff = 24'd14222764;
            12'd1526: coeff = 24'd14232006;
            12'd1527: coeff = 24'd14241234;
            12'd1528: coeff = 24'd14250448;
            12'd1529: coeff = 24'd14259648;
            12'd1530: coeff = 24'd14268834;
            12'd1531: coeff = 24'd14278007;
            12'd1532: coeff = 24'd14287166;
            12'd1533: coeff = 24'd14296310;
            12'd1534: coeff = 24'd14305441;
            12'd1535: coeff = 24'd14314558;
            12'd1536: coeff = 24'd14323661;
            12'd1537: coeff = 24'd14332750;
            12'd1538: coeff = 24'd14341825;
            12'd1539: coeff = 24'd14350886;
            12'd1540: coeff = 24'd14359933;
            12'd1541: coeff = 24'd14368966;
            12'd1542: coeff = 24'd14377985;
            12'd1543: coeff = 24'd14386990;
            12'd1544: coeff = 24'd14395980;
            12'd1545: coeff = 24'd14404957;
            12'd1546: coeff = 24'd14413919;
            12'd1547: coeff = 24'd14422867;
            12'd1548: coeff = 24'd14431801;
            12'd1549: coeff = 24'd14440721;
            12'd1550: coeff = 24'd14449626;
            12'd1551: coeff = 24'd14458517;
            12'd1552: coeff = 24'd14467394;
            12'd1553: coeff = 24'd14476257;
            12'd1554: coeff = 24'd14485105;
            12'd1555: coeff = 24'd14493939;
            12'd1556: coeff = 24'd14502758;
            12'd1557: coeff = 24'd14511564;
            12'd1558: coeff = 24'd14520354;
            12'd1559: coeff = 24'd14529130;
            12'd1560: coeff = 24'd14537892;
            12'd1561: coeff = 24'd14546640;
            12'd1562: coeff = 24'd14555372;
            12'd1563: coeff = 24'd14564091;
            12'd1564: coeff = 24'd14572795;
            12'd1565: coeff = 24'd14581484;
            12'd1566: coeff = 24'd14590158;
            12'd1567: coeff = 24'd14598818;
            12'd1568: coeff = 24'd14607464;
            12'd1569: coeff = 24'd14616095;
            12'd1570: coeff = 24'd14624711;
            12'd1571: coeff = 24'd14633312;
            12'd1572: coeff = 24'd14641899;
            12'd1573: coeff = 24'd14650471;
            12'd1574: coeff = 24'd14659028;
            12'd1575: coeff = 24'd14667571;
            12'd1576: coeff = 24'd14676098;
            12'd1577: coeff = 24'd14684611;
            12'd1578: coeff = 24'd14693110;
            12'd1579: coeff = 24'd14701593;
            12'd1580: coeff = 24'd14710061;
            12'd1581: coeff = 24'd14718515;
            12'd1582: coeff = 24'd14726953;
            12'd1583: coeff = 24'd14735377;
            12'd1584: coeff = 24'd14743786;
            12'd1585: coeff = 24'd14752180;
            12'd1586: coeff = 24'd14760558;
            12'd1587: coeff = 24'd14768922;
            12'd1588: coeff = 24'd14777271;
            12'd1589: coeff = 24'd14785605;
            12'd1590: coeff = 24'd14793923;
            12'd1591: coeff = 24'd14802227;
            12'd1592: coeff = 24'd14810515;
            12'd1593: coeff = 24'd14818789;
            12'd1594: coeff = 24'd14827047;
            12'd1595: coeff = 24'd14835290;
            12'd1596: coeff = 24'd14843518;
            12'd1597: coeff = 24'd14851731;
            12'd1598: coeff = 24'd14859928;
            12'd1599: coeff = 24'd14868111;
            12'd1600: coeff = 24'd14876278;
            12'd1601: coeff = 24'd14884429;
            12'd1602: coeff = 24'd14892566;
            12'd1603: coeff = 24'd14900687;
            12'd1604: coeff = 24'd14908793;
            12'd1605: coeff = 24'd14916883;
            12'd1606: coeff = 24'd14924958;
            12'd1607: coeff = 24'd14933018;
            12'd1608: coeff = 24'd14941062;
            12'd1609: coeff = 24'd14949091;
            12'd1610: coeff = 24'd14957105;
            12'd1611: coeff = 24'd14965102;
            12'd1612: coeff = 24'd14973085;
            12'd1613: coeff = 24'd14981052;
            12'd1614: coeff = 24'd14989003;
            12'd1615: coeff = 24'd14996939;
            12'd1616: coeff = 24'd15004860;
            12'd1617: coeff = 24'd15012764;
            12'd1618: coeff = 24'd15020654;
            12'd1619: coeff = 24'd15028527;
            12'd1620: coeff = 24'd15036385;
            12'd1621: coeff = 24'd15044227;
            12'd1622: coeff = 24'd15052054;
            12'd1623: coeff = 24'd15059865;
            12'd1624: coeff = 24'd15067660;
            12'd1625: coeff = 24'd15075440;
            12'd1626: coeff = 24'd15083203;
            12'd1627: coeff = 24'd15090951;
            12'd1628: coeff = 24'd15098684;
            12'd1629: coeff = 24'd15106400;
            12'd1630: coeff = 24'd15114101;
            12'd1631: coeff = 24'd15121785;
            12'd1632: coeff = 24'd15129454;
            12'd1633: coeff = 24'd15137107;
            12'd1634: coeff = 24'd15144745;
            12'd1635: coeff = 24'd15152366;
            12'd1636: coeff = 24'd15159971;
            12'd1637: coeff = 24'd15167560;
            12'd1638: coeff = 24'd15175134;
            12'd1639: coeff = 24'd15182691;
            12'd1640: coeff = 24'd15190233;
            12'd1641: coeff = 24'd15197758;
            12'd1642: coeff = 24'd15205268;
            12'd1643: coeff = 24'd15212761;
            12'd1644: coeff = 24'd15220238;
            12'd1645: coeff = 24'd15227700;
            12'd1646: coeff = 24'd15235145;
            12'd1647: coeff = 24'd15242574;
            12'd1648: coeff = 24'd15249987;
            12'd1649: coeff = 24'd15257383;
            12'd1650: coeff = 24'd15264764;
            12'd1651: coeff = 24'd15272128;
            12'd1652: coeff = 24'd15279476;
            12'd1653: coeff = 24'd15286808;
            12'd1654: coeff = 24'd15294124;
            12'd1655: coeff = 24'd15301423;
            12'd1656: coeff = 24'd15308707;
            12'd1657: coeff = 24'd15315973;
            12'd1658: coeff = 24'd15323224;
            12'd1659: coeff = 24'd15330458;
            12'd1660: coeff = 24'd15337676;
            12'd1661: coeff = 24'd15344878;
            12'd1662: coeff = 24'd15352063;
            12'd1663: coeff = 24'd15359231;
            12'd1664: coeff = 24'd15366384;
            12'd1665: coeff = 24'd15373520;
            12'd1666: coeff = 24'd15380639;
            12'd1667: coeff = 24'd15387742;
            12'd1668: coeff = 24'd15394829;
            12'd1669: coeff = 24'd15401899;
            12'd1670: coeff = 24'd15408952;
            12'd1671: coeff = 24'd15415989;
            12'd1672: coeff = 24'd15423010;
            12'd1673: coeff = 24'd15430014;
            12'd1674: coeff = 24'd15437001;
            12'd1675: coeff = 24'd15443972;
            12'd1676: coeff = 24'd15450926;
            12'd1677: coeff = 24'd15457863;
            12'd1678: coeff = 24'd15464784;
            12'd1679: coeff = 24'd15471688;
            12'd1680: coeff = 24'd15478576;
            12'd1681: coeff = 24'd15485447;
            12'd1682: coeff = 24'd15492301;
            12'd1683: coeff = 24'd15499138;
            12'd1684: coeff = 24'd15505959;
            12'd1685: coeff = 24'd15512763;
            12'd1686: coeff = 24'd15519550;
            12'd1687: coeff = 24'd15526320;
            12'd1688: coeff = 24'd15533074;
            12'd1689: coeff = 24'd15539810;
            12'd1690: coeff = 24'd15546530;
            12'd1691: coeff = 24'd15553233;
            12'd1692: coeff = 24'd15559919;
            12'd1693: coeff = 24'd15566589;
            12'd1694: coeff = 24'd15573241;
            12'd1695: coeff = 24'd15579876;
            12'd1696: coeff = 24'd15586495;
            12'd1697: coeff = 24'd15593097;
            12'd1698: coeff = 24'd15599681;
            12'd1699: coeff = 24'd15606249;
            12'd1700: coeff = 24'd15612800;
            12'd1701: coeff = 24'd15619333;
            12'd1702: coeff = 24'd15625850;
            12'd1703: coeff = 24'd15632349;
            12'd1704: coeff = 24'd15638832;
            12'd1705: coeff = 24'd15645297;
            12'd1706: coeff = 24'd15651746;
            12'd1707: coeff = 24'd15658177;
            12'd1708: coeff = 24'd15664591;
            12'd1709: coeff = 24'd15670988;
            12'd1710: coeff = 24'd15677368;
            12'd1711: coeff = 24'd15683731;
            12'd1712: coeff = 24'd15690076;
            12'd1713: coeff = 24'd15696405;
            12'd1714: coeff = 24'd15702716;
            12'd1715: coeff = 24'd15709010;
            12'd1716: coeff = 24'd15715287;
            12'd1717: coeff = 24'd15721546;
            12'd1718: coeff = 24'd15727788;
            12'd1719: coeff = 24'd15734013;
            12'd1720: coeff = 24'd15740221;
            12'd1721: coeff = 24'd15746411;
            12'd1722: coeff = 24'd15752584;
            12'd1723: coeff = 24'd15758740;
            12'd1724: coeff = 24'd15764878;
            12'd1725: coeff = 24'd15770999;
            12'd1726: coeff = 24'd15777102;
            12'd1727: coeff = 24'd15783189;
            12'd1728: coeff = 24'd15789257;
            12'd1729: coeff = 24'd15795309;
            12'd1730: coeff = 24'd15801343;
            12'd1731: coeff = 24'd15807359;
            12'd1732: coeff = 24'd15813358;
            12'd1733: coeff = 24'd15819340;
            12'd1734: coeff = 24'd15825304;
            12'd1735: coeff = 24'd15831250;
            12'd1736: coeff = 24'd15837179;
            12'd1737: coeff = 24'd15843090;
            12'd1738: coeff = 24'd15848984;
            12'd1739: coeff = 24'd15854861;
            12'd1740: coeff = 24'd15860719;
            12'd1741: coeff = 24'd15866561;
            12'd1742: coeff = 24'd15872384;
            12'd1743: coeff = 24'd15878190;
            12'd1744: coeff = 24'd15883978;
            12'd1745: coeff = 24'd15889749;
            12'd1746: coeff = 24'd15895502;
            12'd1747: coeff = 24'd15901237;
            12'd1748: coeff = 24'd15906955;
            12'd1749: coeff = 24'd15912655;
            12'd1750: coeff = 24'd15918337;
            12'd1751: coeff = 24'd15924002;
            12'd1752: coeff = 24'd15929648;
            12'd1753: coeff = 24'd15935277;
            12'd1754: coeff = 24'd15940889;
            12'd1755: coeff = 24'd15946482;
            12'd1756: coeff = 24'd15952058;
            12'd1757: coeff = 24'd15957616;
            12'd1758: coeff = 24'd15963156;
            12'd1759: coeff = 24'd15968678;
            12'd1760: coeff = 24'd15974182;
            12'd1761: coeff = 24'd15979669;
            12'd1762: coeff = 24'd15985137;
            12'd1763: coeff = 24'd15990588;
            12'd1764: coeff = 24'd15996021;
            12'd1765: coeff = 24'd16001436;
            12'd1766: coeff = 24'd16006833;
            12'd1767: coeff = 24'd16012212;
            12'd1768: coeff = 24'd16017573;
            12'd1769: coeff = 24'd16022916;
            12'd1770: coeff = 24'd16028242;
            12'd1771: coeff = 24'd16033549;
            12'd1772: coeff = 24'd16038838;
            12'd1773: coeff = 24'd16044109;
            12'd1774: coeff = 24'd16049362;
            12'd1775: coeff = 24'd16054598;
            12'd1776: coeff = 24'd16059815;
            12'd1777: coeff = 24'd16065014;
            12'd1778: coeff = 24'd16070195;
            12'd1779: coeff = 24'd16075358;
            12'd1780: coeff = 24'd16080502;
            12'd1781: coeff = 24'd16085629;
            12'd1782: coeff = 24'd16090738;
            12'd1783: coeff = 24'd16095828;
            12'd1784: coeff = 24'd16100900;
            12'd1785: coeff = 24'd16105954;
            12'd1786: coeff = 24'd16110990;
            12'd1787: coeff = 24'd16116008;
            12'd1788: coeff = 24'd16121008;
            12'd1789: coeff = 24'd16125989;
            12'd1790: coeff = 24'd16130952;
            12'd1791: coeff = 24'd16135897;
            12'd1792: coeff = 24'd16140824;
            12'd1793: coeff = 24'd16145732;
            12'd1794: coeff = 24'd16150623;
            12'd1795: coeff = 24'd16155494;
            12'd1796: coeff = 24'd16160348;
            12'd1797: coeff = 24'd16165183;
            12'd1798: coeff = 24'd16170000;
            12'd1799: coeff = 24'd16174799;
            12'd1800: coeff = 24'd16179580;
            12'd1801: coeff = 24'd16184342;
            12'd1802: coeff = 24'd16189085;
            12'd1803: coeff = 24'd16193811;
            12'd1804: coeff = 24'd16198517;
            12'd1805: coeff = 24'd16203206;
            12'd1806: coeff = 24'd16207876;
            12'd1807: coeff = 24'd16212528;
            12'd1808: coeff = 24'd16217161;
            12'd1809: coeff = 24'd16221776;
            12'd1810: coeff = 24'd16226373;
            12'd1811: coeff = 24'd16230951;
            12'd1812: coeff = 24'd16235510;
            12'd1813: coeff = 24'd16240051;
            12'd1814: coeff = 24'd16244574;
            12'd1815: coeff = 24'd16249078;
            12'd1816: coeff = 24'd16253563;
            12'd1817: coeff = 24'd16258031;
            12'd1818: coeff = 24'd16262479;
            12'd1819: coeff = 24'd16266909;
            12'd1820: coeff = 24'd16271321;
            12'd1821: coeff = 24'd16275713;
            12'd1822: coeff = 24'd16280088;
            12'd1823: coeff = 24'd16284444;
            12'd1824: coeff = 24'd16288781;
            12'd1825: coeff = 24'd16293099;
            12'd1826: coeff = 24'd16297399;
            12'd1827: coeff = 24'd16301681;
            12'd1828: coeff = 24'd16305943;
            12'd1829: coeff = 24'd16310187;
            12'd1830: coeff = 24'd16314413;
            12'd1831: coeff = 24'd16318619;
            12'd1832: coeff = 24'd16322808;
            12'd1833: coeff = 24'd16326977;
            12'd1834: coeff = 24'd16331128;
            12'd1835: coeff = 24'd16335260;
            12'd1836: coeff = 24'd16339373;
            12'd1837: coeff = 24'd16343468;
            12'd1838: coeff = 24'd16347543;
            12'd1839: coeff = 24'd16351601;
            12'd1840: coeff = 24'd16355639;
            12'd1841: coeff = 24'd16359659;
            12'd1842: coeff = 24'd16363659;
            12'd1843: coeff = 24'd16367642;
            12'd1844: coeff = 24'd16371605;
            12'd1845: coeff = 24'd16375549;
            12'd1846: coeff = 24'd16379475;
            12'd1847: coeff = 24'd16383382;
            12'd1848: coeff = 24'd16387270;
            12'd1849: coeff = 24'd16391139;
            12'd1850: coeff = 24'd16394990;
            12'd1851: coeff = 24'd16398821;
            12'd1852: coeff = 24'd16402634;
            12'd1853: coeff = 24'd16406428;
            12'd1854: coeff = 24'd16410203;
            12'd1855: coeff = 24'd16413959;
            12'd1856: coeff = 24'd16417696;
            12'd1857: coeff = 24'd16421414;
            12'd1858: coeff = 24'd16425114;
            12'd1859: coeff = 24'd16428794;
            12'd1860: coeff = 24'd16432455;
            12'd1861: coeff = 24'd16436098;
            12'd1862: coeff = 24'd16439722;
            12'd1863: coeff = 24'd16443326;
            12'd1864: coeff = 24'd16446912;
            12'd1865: coeff = 24'd16450479;
            12'd1866: coeff = 24'd16454027;
            12'd1867: coeff = 24'd16457555;
            12'd1868: coeff = 24'd16461065;
            12'd1869: coeff = 24'd16464556;
            12'd1870: coeff = 24'd16468028;
            12'd1871: coeff = 24'd16471480;
            12'd1872: coeff = 24'd16474914;
            12'd1873: coeff = 24'd16478329;
            12'd1874: coeff = 24'd16481724;
            12'd1875: coeff = 24'd16485101;
            12'd1876: coeff = 24'd16488458;
            12'd1877: coeff = 24'd16491797;
            12'd1878: coeff = 24'd16495116;
            12'd1879: coeff = 24'd16498417;
            12'd1880: coeff = 24'd16501698;
            12'd1881: coeff = 24'd16504960;
            12'd1882: coeff = 24'd16508203;
            12'd1883: coeff = 24'd16511427;
            12'd1884: coeff = 24'd16514631;
            12'd1885: coeff = 24'd16517817;
            12'd1886: coeff = 24'd16520983;
            12'd1887: coeff = 24'd16524131;
            12'd1888: coeff = 24'd16527259;
            12'd1889: coeff = 24'd16530368;
            12'd1890: coeff = 24'd16533458;
            12'd1891: coeff = 24'd16536528;
            12'd1892: coeff = 24'd16539580;
            12'd1893: coeff = 24'd16542612;
            12'd1894: coeff = 24'd16545625;
            12'd1895: coeff = 24'd16548619;
            12'd1896: coeff = 24'd16551594;
            12'd1897: coeff = 24'd16554549;
            12'd1898: coeff = 24'd16557486;
            12'd1899: coeff = 24'd16560403;
            12'd1900: coeff = 24'd16563300;
            12'd1901: coeff = 24'd16566179;
            12'd1902: coeff = 24'd16569038;
            12'd1903: coeff = 24'd16571878;
            12'd1904: coeff = 24'd16574699;
            12'd1905: coeff = 24'd16577500;
            12'd1906: coeff = 24'd16580283;
            12'd1907: coeff = 24'd16583046;
            12'd1908: coeff = 24'd16585789;
            12'd1909: coeff = 24'd16588514;
            12'd1910: coeff = 24'd16591219;
            12'd1911: coeff = 24'd16593904;
            12'd1912: coeff = 24'd16596571;
            12'd1913: coeff = 24'd16599218;
            12'd1914: coeff = 24'd16601845;
            12'd1915: coeff = 24'd16604454;
            12'd1916: coeff = 24'd16607043;
            12'd1917: coeff = 24'd16609613;
            12'd1918: coeff = 24'd16612163;
            12'd1919: coeff = 24'd16614694;
            12'd1920: coeff = 24'd16617206;
            12'd1921: coeff = 24'd16619698;
            12'd1922: coeff = 24'd16622171;
            12'd1923: coeff = 24'd16624624;
            12'd1924: coeff = 24'd16627058;
            12'd1925: coeff = 24'd16629473;
            12'd1926: coeff = 24'd16631868;
            12'd1927: coeff = 24'd16634244;
            12'd1928: coeff = 24'd16636601;
            12'd1929: coeff = 24'd16638938;
            12'd1930: coeff = 24'd16641256;
            12'd1931: coeff = 24'd16643554;
            12'd1932: coeff = 24'd16645833;
            12'd1933: coeff = 24'd16648092;
            12'd1934: coeff = 24'd16650332;
            12'd1935: coeff = 24'd16652552;
            12'd1936: coeff = 24'd16654753;
            12'd1937: coeff = 24'd16656935;
            12'd1938: coeff = 24'd16659097;
            12'd1939: coeff = 24'd16661240;
            12'd1940: coeff = 24'd16663363;
            12'd1941: coeff = 24'd16665466;
            12'd1942: coeff = 24'd16667550;
            12'd1943: coeff = 24'd16669615;
            12'd1944: coeff = 24'd16671660;
            12'd1945: coeff = 24'd16673686;
            12'd1946: coeff = 24'd16675692;
            12'd1947: coeff = 24'd16677679;
            12'd1948: coeff = 24'd16679646;
            12'd1949: coeff = 24'd16681594;
            12'd1950: coeff = 24'd16683522;
            12'd1951: coeff = 24'd16685430;
            12'd1952: coeff = 24'd16687319;
            12'd1953: coeff = 24'd16689189;
            12'd1954: coeff = 24'd16691039;
            12'd1955: coeff = 24'd16692869;
            12'd1956: coeff = 24'd16694680;
            12'd1957: coeff = 24'd16696471;
            12'd1958: coeff = 24'd16698243;
            12'd1959: coeff = 24'd16699995;
            12'd1960: coeff = 24'd16701728;
            12'd1961: coeff = 24'd16703441;
            12'd1962: coeff = 24'd16705134;
            12'd1963: coeff = 24'd16706808;
            12'd1964: coeff = 24'd16708463;
            12'd1965: coeff = 24'd16710097;
            12'd1966: coeff = 24'd16711713;
            12'd1967: coeff = 24'd16713308;
            12'd1968: coeff = 24'd16714884;
            12'd1969: coeff = 24'd16716440;
            12'd1970: coeff = 24'd16717977;
            12'd1971: coeff = 24'd16719494;
            12'd1972: coeff = 24'd16720992;
            12'd1973: coeff = 24'd16722470;
            12'd1974: coeff = 24'd16723928;
            12'd1975: coeff = 24'd16725367;
            12'd1976: coeff = 24'd16726786;
            12'd1977: coeff = 24'd16728185;
            12'd1978: coeff = 24'd16729565;
            12'd1979: coeff = 24'd16730925;
            12'd1980: coeff = 24'd16732265;
            12'd1981: coeff = 24'd16733586;
            12'd1982: coeff = 24'd16734887;
            12'd1983: coeff = 24'd16736169;
            12'd1984: coeff = 24'd16737431;
            12'd1985: coeff = 24'd16738673;
            12'd1986: coeff = 24'd16739896;
            12'd1987: coeff = 24'd16741099;
            12'd1988: coeff = 24'd16742282;
            12'd1989: coeff = 24'd16743445;
            12'd1990: coeff = 24'd16744589;
            12'd1991: coeff = 24'd16745714;
            12'd1992: coeff = 24'd16746818;
            12'd1993: coeff = 24'd16747903;
            12'd1994: coeff = 24'd16748968;
            12'd1995: coeff = 24'd16750014;
            12'd1996: coeff = 24'd16751040;
            12'd1997: coeff = 24'd16752046;
            12'd1998: coeff = 24'd16753032;
            12'd1999: coeff = 24'd16753999;
            12'd2000: coeff = 24'd16754946;
            12'd2001: coeff = 24'd16755874;
            12'd2002: coeff = 24'd16756781;
            12'd2003: coeff = 24'd16757669;
            12'd2004: coeff = 24'd16758538;
            12'd2005: coeff = 24'd16759386;
            12'd2006: coeff = 24'd16760215;
            12'd2007: coeff = 24'd16761024;
            12'd2008: coeff = 24'd16761814;
            12'd2009: coeff = 24'd16762583;
            12'd2010: coeff = 24'd16763333;
            12'd2011: coeff = 24'd16764064;
            12'd2012: coeff = 24'd16764774;
            12'd2013: coeff = 24'd16765465;
            12'd2014: coeff = 24'd16766136;
            12'd2015: coeff = 24'd16766788;
            12'd2016: coeff = 24'd16767420;
            12'd2017: coeff = 24'd16768031;
            12'd2018: coeff = 24'd16768624;
            12'd2019: coeff = 24'd16769196;
            12'd2020: coeff = 24'd16769749;
            12'd2021: coeff = 24'd16770282;
            12'd2022: coeff = 24'd16770795;
            12'd2023: coeff = 24'd16771289;
            12'd2024: coeff = 24'd16771763;
            12'd2025: coeff = 24'd16772217;
            12'd2026: coeff = 24'd16772651;
            12'd2027: coeff = 24'd16773066;
            12'd2028: coeff = 24'd16773461;
            12'd2029: coeff = 24'd16773836;
            12'd2030: coeff = 24'd16774192;
            12'd2031: coeff = 24'd16774527;
            12'd2032: coeff = 24'd16774843;
            12'd2033: coeff = 24'd16775139;
            12'd2034: coeff = 24'd16775416;
            12'd2035: coeff = 24'd16775673;
            12'd2036: coeff = 24'd16775910;
            12'd2037: coeff = 24'd16776127;
            12'd2038: coeff = 24'd16776324;
            12'd2039: coeff = 24'd16776502;
            12'd2040: coeff = 24'd16776660;
            12'd2041: coeff = 24'd16776798;
            12'd2042: coeff = 24'd16776917;
            12'd2043: coeff = 24'd16777016;
            12'd2044: coeff = 24'd16777095;
            12'd2045: coeff = 24'd16777154;
            12'd2046: coeff = 24'd16777193;
            12'd2047: coeff = 24'd16777213;
            12'd2048: coeff = 24'd16777213;
            12'd2049: coeff = 24'd16777193;
            12'd2050: coeff = 24'd16777154;
            12'd2051: coeff = 24'd16777095;
            12'd2052: coeff = 24'd16777016;
            12'd2053: coeff = 24'd16776917;
            12'd2054: coeff = 24'd16776798;
            12'd2055: coeff = 24'd16776660;
            12'd2056: coeff = 24'd16776502;
            12'd2057: coeff = 24'd16776324;
            12'd2058: coeff = 24'd16776127;
            12'd2059: coeff = 24'd16775910;
            12'd2060: coeff = 24'd16775673;
            12'd2061: coeff = 24'd16775416;
            12'd2062: coeff = 24'd16775139;
            12'd2063: coeff = 24'd16774843;
            12'd2064: coeff = 24'd16774527;
            12'd2065: coeff = 24'd16774192;
            12'd2066: coeff = 24'd16773836;
            12'd2067: coeff = 24'd16773461;
            12'd2068: coeff = 24'd16773066;
            12'd2069: coeff = 24'd16772651;
            12'd2070: coeff = 24'd16772217;
            12'd2071: coeff = 24'd16771763;
            12'd2072: coeff = 24'd16771289;
            12'd2073: coeff = 24'd16770795;
            12'd2074: coeff = 24'd16770282;
            12'd2075: coeff = 24'd16769749;
            12'd2076: coeff = 24'd16769196;
            12'd2077: coeff = 24'd16768624;
            12'd2078: coeff = 24'd16768031;
            12'd2079: coeff = 24'd16767420;
            12'd2080: coeff = 24'd16766788;
            12'd2081: coeff = 24'd16766136;
            12'd2082: coeff = 24'd16765465;
            12'd2083: coeff = 24'd16764774;
            12'd2084: coeff = 24'd16764064;
            12'd2085: coeff = 24'd16763333;
            12'd2086: coeff = 24'd16762583;
            12'd2087: coeff = 24'd16761814;
            12'd2088: coeff = 24'd16761024;
            12'd2089: coeff = 24'd16760215;
            12'd2090: coeff = 24'd16759386;
            12'd2091: coeff = 24'd16758538;
            12'd2092: coeff = 24'd16757669;
            12'd2093: coeff = 24'd16756781;
            12'd2094: coeff = 24'd16755874;
            12'd2095: coeff = 24'd16754946;
            12'd2096: coeff = 24'd16753999;
            12'd2097: coeff = 24'd16753032;
            12'd2098: coeff = 24'd16752046;
            12'd2099: coeff = 24'd16751040;
            12'd2100: coeff = 24'd16750014;
            12'd2101: coeff = 24'd16748968;
            12'd2102: coeff = 24'd16747903;
            12'd2103: coeff = 24'd16746818;
            12'd2104: coeff = 24'd16745714;
            12'd2105: coeff = 24'd16744589;
            12'd2106: coeff = 24'd16743445;
            12'd2107: coeff = 24'd16742282;
            12'd2108: coeff = 24'd16741099;
            12'd2109: coeff = 24'd16739896;
            12'd2110: coeff = 24'd16738673;
            12'd2111: coeff = 24'd16737431;
            12'd2112: coeff = 24'd16736169;
            12'd2113: coeff = 24'd16734887;
            12'd2114: coeff = 24'd16733586;
            12'd2115: coeff = 24'd16732265;
            12'd2116: coeff = 24'd16730925;
            12'd2117: coeff = 24'd16729565;
            12'd2118: coeff = 24'd16728185;
            12'd2119: coeff = 24'd16726786;
            12'd2120: coeff = 24'd16725367;
            12'd2121: coeff = 24'd16723928;
            12'd2122: coeff = 24'd16722470;
            12'd2123: coeff = 24'd16720992;
            12'd2124: coeff = 24'd16719494;
            12'd2125: coeff = 24'd16717977;
            12'd2126: coeff = 24'd16716440;
            12'd2127: coeff = 24'd16714884;
            12'd2128: coeff = 24'd16713308;
            12'd2129: coeff = 24'd16711713;
            12'd2130: coeff = 24'd16710097;
            12'd2131: coeff = 24'd16708463;
            12'd2132: coeff = 24'd16706808;
            12'd2133: coeff = 24'd16705134;
            12'd2134: coeff = 24'd16703441;
            12'd2135: coeff = 24'd16701728;
            12'd2136: coeff = 24'd16699995;
            12'd2137: coeff = 24'd16698243;
            12'd2138: coeff = 24'd16696471;
            12'd2139: coeff = 24'd16694680;
            12'd2140: coeff = 24'd16692869;
            12'd2141: coeff = 24'd16691039;
            12'd2142: coeff = 24'd16689189;
            12'd2143: coeff = 24'd16687319;
            12'd2144: coeff = 24'd16685430;
            12'd2145: coeff = 24'd16683522;
            12'd2146: coeff = 24'd16681594;
            12'd2147: coeff = 24'd16679646;
            12'd2148: coeff = 24'd16677679;
            12'd2149: coeff = 24'd16675692;
            12'd2150: coeff = 24'd16673686;
            12'd2151: coeff = 24'd16671660;
            12'd2152: coeff = 24'd16669615;
            12'd2153: coeff = 24'd16667550;
            12'd2154: coeff = 24'd16665466;
            12'd2155: coeff = 24'd16663363;
            12'd2156: coeff = 24'd16661240;
            12'd2157: coeff = 24'd16659097;
            12'd2158: coeff = 24'd16656935;
            12'd2159: coeff = 24'd16654753;
            12'd2160: coeff = 24'd16652552;
            12'd2161: coeff = 24'd16650332;
            12'd2162: coeff = 24'd16648092;
            12'd2163: coeff = 24'd16645833;
            12'd2164: coeff = 24'd16643554;
            12'd2165: coeff = 24'd16641256;
            12'd2166: coeff = 24'd16638938;
            12'd2167: coeff = 24'd16636601;
            12'd2168: coeff = 24'd16634244;
            12'd2169: coeff = 24'd16631868;
            12'd2170: coeff = 24'd16629473;
            12'd2171: coeff = 24'd16627058;
            12'd2172: coeff = 24'd16624624;
            12'd2173: coeff = 24'd16622171;
            12'd2174: coeff = 24'd16619698;
            12'd2175: coeff = 24'd16617206;
            12'd2176: coeff = 24'd16614694;
            12'd2177: coeff = 24'd16612163;
            12'd2178: coeff = 24'd16609613;
            12'd2179: coeff = 24'd16607043;
            12'd2180: coeff = 24'd16604454;
            12'd2181: coeff = 24'd16601845;
            12'd2182: coeff = 24'd16599218;
            12'd2183: coeff = 24'd16596571;
            12'd2184: coeff = 24'd16593904;
            12'd2185: coeff = 24'd16591219;
            12'd2186: coeff = 24'd16588514;
            12'd2187: coeff = 24'd16585789;
            12'd2188: coeff = 24'd16583046;
            12'd2189: coeff = 24'd16580283;
            12'd2190: coeff = 24'd16577500;
            12'd2191: coeff = 24'd16574699;
            12'd2192: coeff = 24'd16571878;
            12'd2193: coeff = 24'd16569038;
            12'd2194: coeff = 24'd16566179;
            12'd2195: coeff = 24'd16563300;
            12'd2196: coeff = 24'd16560403;
            12'd2197: coeff = 24'd16557486;
            12'd2198: coeff = 24'd16554549;
            12'd2199: coeff = 24'd16551594;
            12'd2200: coeff = 24'd16548619;
            12'd2201: coeff = 24'd16545625;
            12'd2202: coeff = 24'd16542612;
            12'd2203: coeff = 24'd16539580;
            12'd2204: coeff = 24'd16536528;
            12'd2205: coeff = 24'd16533458;
            12'd2206: coeff = 24'd16530368;
            12'd2207: coeff = 24'd16527259;
            12'd2208: coeff = 24'd16524131;
            12'd2209: coeff = 24'd16520983;
            12'd2210: coeff = 24'd16517817;
            12'd2211: coeff = 24'd16514631;
            12'd2212: coeff = 24'd16511427;
            12'd2213: coeff = 24'd16508203;
            12'd2214: coeff = 24'd16504960;
            12'd2215: coeff = 24'd16501698;
            12'd2216: coeff = 24'd16498417;
            12'd2217: coeff = 24'd16495116;
            12'd2218: coeff = 24'd16491797;
            12'd2219: coeff = 24'd16488458;
            12'd2220: coeff = 24'd16485101;
            12'd2221: coeff = 24'd16481724;
            12'd2222: coeff = 24'd16478329;
            12'd2223: coeff = 24'd16474914;
            12'd2224: coeff = 24'd16471480;
            12'd2225: coeff = 24'd16468028;
            12'd2226: coeff = 24'd16464556;
            12'd2227: coeff = 24'd16461065;
            12'd2228: coeff = 24'd16457555;
            12'd2229: coeff = 24'd16454027;
            12'd2230: coeff = 24'd16450479;
            12'd2231: coeff = 24'd16446912;
            12'd2232: coeff = 24'd16443326;
            12'd2233: coeff = 24'd16439722;
            12'd2234: coeff = 24'd16436098;
            12'd2235: coeff = 24'd16432455;
            12'd2236: coeff = 24'd16428794;
            12'd2237: coeff = 24'd16425114;
            12'd2238: coeff = 24'd16421414;
            12'd2239: coeff = 24'd16417696;
            12'd2240: coeff = 24'd16413959;
            12'd2241: coeff = 24'd16410203;
            12'd2242: coeff = 24'd16406428;
            12'd2243: coeff = 24'd16402634;
            12'd2244: coeff = 24'd16398821;
            12'd2245: coeff = 24'd16394990;
            12'd2246: coeff = 24'd16391139;
            12'd2247: coeff = 24'd16387270;
            12'd2248: coeff = 24'd16383382;
            12'd2249: coeff = 24'd16379475;
            12'd2250: coeff = 24'd16375549;
            12'd2251: coeff = 24'd16371605;
            12'd2252: coeff = 24'd16367642;
            12'd2253: coeff = 24'd16363659;
            12'd2254: coeff = 24'd16359659;
            12'd2255: coeff = 24'd16355639;
            12'd2256: coeff = 24'd16351601;
            12'd2257: coeff = 24'd16347543;
            12'd2258: coeff = 24'd16343468;
            12'd2259: coeff = 24'd16339373;
            12'd2260: coeff = 24'd16335260;
            12'd2261: coeff = 24'd16331128;
            12'd2262: coeff = 24'd16326977;
            12'd2263: coeff = 24'd16322808;
            12'd2264: coeff = 24'd16318619;
            12'd2265: coeff = 24'd16314413;
            12'd2266: coeff = 24'd16310187;
            12'd2267: coeff = 24'd16305943;
            12'd2268: coeff = 24'd16301681;
            12'd2269: coeff = 24'd16297399;
            12'd2270: coeff = 24'd16293099;
            12'd2271: coeff = 24'd16288781;
            12'd2272: coeff = 24'd16284444;
            12'd2273: coeff = 24'd16280088;
            12'd2274: coeff = 24'd16275713;
            12'd2275: coeff = 24'd16271321;
            12'd2276: coeff = 24'd16266909;
            12'd2277: coeff = 24'd16262479;
            12'd2278: coeff = 24'd16258031;
            12'd2279: coeff = 24'd16253563;
            12'd2280: coeff = 24'd16249078;
            12'd2281: coeff = 24'd16244574;
            12'd2282: coeff = 24'd16240051;
            12'd2283: coeff = 24'd16235510;
            12'd2284: coeff = 24'd16230951;
            12'd2285: coeff = 24'd16226373;
            12'd2286: coeff = 24'd16221776;
            12'd2287: coeff = 24'd16217161;
            12'd2288: coeff = 24'd16212528;
            12'd2289: coeff = 24'd16207876;
            12'd2290: coeff = 24'd16203206;
            12'd2291: coeff = 24'd16198517;
            12'd2292: coeff = 24'd16193811;
            12'd2293: coeff = 24'd16189085;
            12'd2294: coeff = 24'd16184342;
            12'd2295: coeff = 24'd16179580;
            12'd2296: coeff = 24'd16174799;
            12'd2297: coeff = 24'd16170000;
            12'd2298: coeff = 24'd16165183;
            12'd2299: coeff = 24'd16160348;
            12'd2300: coeff = 24'd16155494;
            12'd2301: coeff = 24'd16150623;
            12'd2302: coeff = 24'd16145732;
            12'd2303: coeff = 24'd16140824;
            12'd2304: coeff = 24'd16135897;
            12'd2305: coeff = 24'd16130952;
            12'd2306: coeff = 24'd16125989;
            12'd2307: coeff = 24'd16121008;
            12'd2308: coeff = 24'd16116008;
            12'd2309: coeff = 24'd16110990;
            12'd2310: coeff = 24'd16105954;
            12'd2311: coeff = 24'd16100900;
            12'd2312: coeff = 24'd16095828;
            12'd2313: coeff = 24'd16090738;
            12'd2314: coeff = 24'd16085629;
            12'd2315: coeff = 24'd16080502;
            12'd2316: coeff = 24'd16075358;
            12'd2317: coeff = 24'd16070195;
            12'd2318: coeff = 24'd16065014;
            12'd2319: coeff = 24'd16059815;
            12'd2320: coeff = 24'd16054598;
            12'd2321: coeff = 24'd16049362;
            12'd2322: coeff = 24'd16044109;
            12'd2323: coeff = 24'd16038838;
            12'd2324: coeff = 24'd16033549;
            12'd2325: coeff = 24'd16028242;
            12'd2326: coeff = 24'd16022916;
            12'd2327: coeff = 24'd16017573;
            12'd2328: coeff = 24'd16012212;
            12'd2329: coeff = 24'd16006833;
            12'd2330: coeff = 24'd16001436;
            12'd2331: coeff = 24'd15996021;
            12'd2332: coeff = 24'd15990588;
            12'd2333: coeff = 24'd15985137;
            12'd2334: coeff = 24'd15979669;
            12'd2335: coeff = 24'd15974182;
            12'd2336: coeff = 24'd15968678;
            12'd2337: coeff = 24'd15963156;
            12'd2338: coeff = 24'd15957616;
            12'd2339: coeff = 24'd15952058;
            12'd2340: coeff = 24'd15946482;
            12'd2341: coeff = 24'd15940889;
            12'd2342: coeff = 24'd15935277;
            12'd2343: coeff = 24'd15929648;
            12'd2344: coeff = 24'd15924002;
            12'd2345: coeff = 24'd15918337;
            12'd2346: coeff = 24'd15912655;
            12'd2347: coeff = 24'd15906955;
            12'd2348: coeff = 24'd15901237;
            12'd2349: coeff = 24'd15895502;
            12'd2350: coeff = 24'd15889749;
            12'd2351: coeff = 24'd15883978;
            12'd2352: coeff = 24'd15878190;
            12'd2353: coeff = 24'd15872384;
            12'd2354: coeff = 24'd15866561;
            12'd2355: coeff = 24'd15860719;
            12'd2356: coeff = 24'd15854861;
            12'd2357: coeff = 24'd15848984;
            12'd2358: coeff = 24'd15843090;
            12'd2359: coeff = 24'd15837179;
            12'd2360: coeff = 24'd15831250;
            12'd2361: coeff = 24'd15825304;
            12'd2362: coeff = 24'd15819340;
            12'd2363: coeff = 24'd15813358;
            12'd2364: coeff = 24'd15807359;
            12'd2365: coeff = 24'd15801343;
            12'd2366: coeff = 24'd15795309;
            12'd2367: coeff = 24'd15789257;
            12'd2368: coeff = 24'd15783189;
            12'd2369: coeff = 24'd15777102;
            12'd2370: coeff = 24'd15770999;
            12'd2371: coeff = 24'd15764878;
            12'd2372: coeff = 24'd15758740;
            12'd2373: coeff = 24'd15752584;
            12'd2374: coeff = 24'd15746411;
            12'd2375: coeff = 24'd15740221;
            12'd2376: coeff = 24'd15734013;
            12'd2377: coeff = 24'd15727788;
            12'd2378: coeff = 24'd15721546;
            12'd2379: coeff = 24'd15715287;
            12'd2380: coeff = 24'd15709010;
            12'd2381: coeff = 24'd15702716;
            12'd2382: coeff = 24'd15696405;
            12'd2383: coeff = 24'd15690076;
            12'd2384: coeff = 24'd15683731;
            12'd2385: coeff = 24'd15677368;
            12'd2386: coeff = 24'd15670988;
            12'd2387: coeff = 24'd15664591;
            12'd2388: coeff = 24'd15658177;
            12'd2389: coeff = 24'd15651746;
            12'd2390: coeff = 24'd15645297;
            12'd2391: coeff = 24'd15638832;
            12'd2392: coeff = 24'd15632349;
            12'd2393: coeff = 24'd15625850;
            12'd2394: coeff = 24'd15619333;
            12'd2395: coeff = 24'd15612800;
            12'd2396: coeff = 24'd15606249;
            12'd2397: coeff = 24'd15599681;
            12'd2398: coeff = 24'd15593097;
            12'd2399: coeff = 24'd15586495;
            12'd2400: coeff = 24'd15579876;
            12'd2401: coeff = 24'd15573241;
            12'd2402: coeff = 24'd15566589;
            12'd2403: coeff = 24'd15559919;
            12'd2404: coeff = 24'd15553233;
            12'd2405: coeff = 24'd15546530;
            12'd2406: coeff = 24'd15539810;
            12'd2407: coeff = 24'd15533074;
            12'd2408: coeff = 24'd15526320;
            12'd2409: coeff = 24'd15519550;
            12'd2410: coeff = 24'd15512763;
            12'd2411: coeff = 24'd15505959;
            12'd2412: coeff = 24'd15499138;
            12'd2413: coeff = 24'd15492301;
            12'd2414: coeff = 24'd15485447;
            12'd2415: coeff = 24'd15478576;
            12'd2416: coeff = 24'd15471688;
            12'd2417: coeff = 24'd15464784;
            12'd2418: coeff = 24'd15457863;
            12'd2419: coeff = 24'd15450926;
            12'd2420: coeff = 24'd15443972;
            12'd2421: coeff = 24'd15437001;
            12'd2422: coeff = 24'd15430014;
            12'd2423: coeff = 24'd15423010;
            12'd2424: coeff = 24'd15415989;
            12'd2425: coeff = 24'd15408952;
            12'd2426: coeff = 24'd15401899;
            12'd2427: coeff = 24'd15394829;
            12'd2428: coeff = 24'd15387742;
            12'd2429: coeff = 24'd15380639;
            12'd2430: coeff = 24'd15373520;
            12'd2431: coeff = 24'd15366384;
            12'd2432: coeff = 24'd15359231;
            12'd2433: coeff = 24'd15352063;
            12'd2434: coeff = 24'd15344878;
            12'd2435: coeff = 24'd15337676;
            12'd2436: coeff = 24'd15330458;
            12'd2437: coeff = 24'd15323224;
            12'd2438: coeff = 24'd15315973;
            12'd2439: coeff = 24'd15308707;
            12'd2440: coeff = 24'd15301423;
            12'd2441: coeff = 24'd15294124;
            12'd2442: coeff = 24'd15286808;
            12'd2443: coeff = 24'd15279476;
            12'd2444: coeff = 24'd15272128;
            12'd2445: coeff = 24'd15264764;
            12'd2446: coeff = 24'd15257383;
            12'd2447: coeff = 24'd15249987;
            12'd2448: coeff = 24'd15242574;
            12'd2449: coeff = 24'd15235145;
            12'd2450: coeff = 24'd15227700;
            12'd2451: coeff = 24'd15220238;
            12'd2452: coeff = 24'd15212761;
            12'd2453: coeff = 24'd15205268;
            12'd2454: coeff = 24'd15197758;
            12'd2455: coeff = 24'd15190233;
            12'd2456: coeff = 24'd15182691;
            12'd2457: coeff = 24'd15175134;
            12'd2458: coeff = 24'd15167560;
            12'd2459: coeff = 24'd15159971;
            12'd2460: coeff = 24'd15152366;
            12'd2461: coeff = 24'd15144745;
            12'd2462: coeff = 24'd15137107;
            12'd2463: coeff = 24'd15129454;
            12'd2464: coeff = 24'd15121785;
            12'd2465: coeff = 24'd15114101;
            12'd2466: coeff = 24'd15106400;
            12'd2467: coeff = 24'd15098684;
            12'd2468: coeff = 24'd15090951;
            12'd2469: coeff = 24'd15083203;
            12'd2470: coeff = 24'd15075440;
            12'd2471: coeff = 24'd15067660;
            12'd2472: coeff = 24'd15059865;
            12'd2473: coeff = 24'd15052054;
            12'd2474: coeff = 24'd15044227;
            12'd2475: coeff = 24'd15036385;
            12'd2476: coeff = 24'd15028527;
            12'd2477: coeff = 24'd15020654;
            12'd2478: coeff = 24'd15012764;
            12'd2479: coeff = 24'd15004860;
            12'd2480: coeff = 24'd14996939;
            12'd2481: coeff = 24'd14989003;
            12'd2482: coeff = 24'd14981052;
            12'd2483: coeff = 24'd14973085;
            12'd2484: coeff = 24'd14965102;
            12'd2485: coeff = 24'd14957105;
            12'd2486: coeff = 24'd14949091;
            12'd2487: coeff = 24'd14941062;
            12'd2488: coeff = 24'd14933018;
            12'd2489: coeff = 24'd14924958;
            12'd2490: coeff = 24'd14916883;
            12'd2491: coeff = 24'd14908793;
            12'd2492: coeff = 24'd14900687;
            12'd2493: coeff = 24'd14892566;
            12'd2494: coeff = 24'd14884429;
            12'd2495: coeff = 24'd14876278;
            12'd2496: coeff = 24'd14868111;
            12'd2497: coeff = 24'd14859928;
            12'd2498: coeff = 24'd14851731;
            12'd2499: coeff = 24'd14843518;
            12'd2500: coeff = 24'd14835290;
            12'd2501: coeff = 24'd14827047;
            12'd2502: coeff = 24'd14818789;
            12'd2503: coeff = 24'd14810515;
            12'd2504: coeff = 24'd14802227;
            12'd2505: coeff = 24'd14793923;
            12'd2506: coeff = 24'd14785605;
            12'd2507: coeff = 24'd14777271;
            12'd2508: coeff = 24'd14768922;
            12'd2509: coeff = 24'd14760558;
            12'd2510: coeff = 24'd14752180;
            12'd2511: coeff = 24'd14743786;
            12'd2512: coeff = 24'd14735377;
            12'd2513: coeff = 24'd14726953;
            12'd2514: coeff = 24'd14718515;
            12'd2515: coeff = 24'd14710061;
            12'd2516: coeff = 24'd14701593;
            12'd2517: coeff = 24'd14693110;
            12'd2518: coeff = 24'd14684611;
            12'd2519: coeff = 24'd14676098;
            12'd2520: coeff = 24'd14667571;
            12'd2521: coeff = 24'd14659028;
            12'd2522: coeff = 24'd14650471;
            12'd2523: coeff = 24'd14641899;
            12'd2524: coeff = 24'd14633312;
            12'd2525: coeff = 24'd14624711;
            12'd2526: coeff = 24'd14616095;
            12'd2527: coeff = 24'd14607464;
            12'd2528: coeff = 24'd14598818;
            12'd2529: coeff = 24'd14590158;
            12'd2530: coeff = 24'd14581484;
            12'd2531: coeff = 24'd14572795;
            12'd2532: coeff = 24'd14564091;
            12'd2533: coeff = 24'd14555372;
            12'd2534: coeff = 24'd14546640;
            12'd2535: coeff = 24'd14537892;
            12'd2536: coeff = 24'd14529130;
            12'd2537: coeff = 24'd14520354;
            12'd2538: coeff = 24'd14511564;
            12'd2539: coeff = 24'd14502758;
            12'd2540: coeff = 24'd14493939;
            12'd2541: coeff = 24'd14485105;
            12'd2542: coeff = 24'd14476257;
            12'd2543: coeff = 24'd14467394;
            12'd2544: coeff = 24'd14458517;
            12'd2545: coeff = 24'd14449626;
            12'd2546: coeff = 24'd14440721;
            12'd2547: coeff = 24'd14431801;
            12'd2548: coeff = 24'd14422867;
            12'd2549: coeff = 24'd14413919;
            12'd2550: coeff = 24'd14404957;
            12'd2551: coeff = 24'd14395980;
            12'd2552: coeff = 24'd14386990;
            12'd2553: coeff = 24'd14377985;
            12'd2554: coeff = 24'd14368966;
            12'd2555: coeff = 24'd14359933;
            12'd2556: coeff = 24'd14350886;
            12'd2557: coeff = 24'd14341825;
            12'd2558: coeff = 24'd14332750;
            12'd2559: coeff = 24'd14323661;
            12'd2560: coeff = 24'd14314558;
            12'd2561: coeff = 24'd14305441;
            12'd2562: coeff = 24'd14296310;
            12'd2563: coeff = 24'd14287166;
            12'd2564: coeff = 24'd14278007;
            12'd2565: coeff = 24'd14268834;
            12'd2566: coeff = 24'd14259648;
            12'd2567: coeff = 24'd14250448;
            12'd2568: coeff = 24'd14241234;
            12'd2569: coeff = 24'd14232006;
            12'd2570: coeff = 24'd14222764;
            12'd2571: coeff = 24'd14213509;
            12'd2572: coeff = 24'd14204240;
            12'd2573: coeff = 24'd14194958;
            12'd2574: coeff = 24'd14185661;
            12'd2575: coeff = 24'd14176351;
            12'd2576: coeff = 24'd14167028;
            12'd2577: coeff = 24'd14157690;
            12'd2578: coeff = 24'd14148340;
            12'd2579: coeff = 24'd14138975;
            12'd2580: coeff = 24'd14129597;
            12'd2581: coeff = 24'd14120206;
            12'd2582: coeff = 24'd14110801;
            12'd2583: coeff = 24'd14101383;
            12'd2584: coeff = 24'd14091951;
            12'd2585: coeff = 24'd14082505;
            12'd2586: coeff = 24'd14073047;
            12'd2587: coeff = 24'd14063575;
            12'd2588: coeff = 24'd14054089;
            12'd2589: coeff = 24'd14044591;
            12'd2590: coeff = 24'd14035079;
            12'd2591: coeff = 24'd14025553;
            12'd2592: coeff = 24'd14016015;
            12'd2593: coeff = 24'd14006463;
            12'd2594: coeff = 24'd13996898;
            12'd2595: coeff = 24'd13987319;
            12'd2596: coeff = 24'd13977728;
            12'd2597: coeff = 24'd13968123;
            12'd2598: coeff = 24'd13958505;
            12'd2599: coeff = 24'd13948875;
            12'd2600: coeff = 24'd13939231;
            12'd2601: coeff = 24'd13929574;
            12'd2602: coeff = 24'd13919903;
            12'd2603: coeff = 24'd13910220;
            12'd2604: coeff = 24'd13900524;
            12'd2605: coeff = 24'd13890815;
            12'd2606: coeff = 24'd13881093;
            12'd2607: coeff = 24'd13871358;
            12'd2608: coeff = 24'd13861610;
            12'd2609: coeff = 24'd13851850;
            12'd2610: coeff = 24'd13842076;
            12'd2611: coeff = 24'd13832289;
            12'd2612: coeff = 24'd13822490;
            12'd2613: coeff = 24'd13812678;
            12'd2614: coeff = 24'd13802853;
            12'd2615: coeff = 24'd13793016;
            12'd2616: coeff = 24'd13783165;
            12'd2617: coeff = 24'd13773302;
            12'd2618: coeff = 24'd13763427;
            12'd2619: coeff = 24'd13753538;
            12'd2620: coeff = 24'd13743637;
            12'd2621: coeff = 24'd13733724;
            12'd2622: coeff = 24'd13723798;
            12'd2623: coeff = 24'd13713859;
            12'd2624: coeff = 24'd13703908;
            12'd2625: coeff = 24'd13693944;
            12'd2626: coeff = 24'd13683968;
            12'd2627: coeff = 24'd13673979;
            12'd2628: coeff = 24'd13663978;
            12'd2629: coeff = 24'd13653964;
            12'd2630: coeff = 24'd13643938;
            12'd2631: coeff = 24'd13633900;
            12'd2632: coeff = 24'd13623849;
            12'd2633: coeff = 24'd13613786;
            12'd2634: coeff = 24'd13603711;
            12'd2635: coeff = 24'd13593623;
            12'd2636: coeff = 24'd13583523;
            12'd2637: coeff = 24'd13573411;
            12'd2638: coeff = 24'd13563287;
            12'd2639: coeff = 24'd13553150;
            12'd2640: coeff = 24'd13543002;
            12'd2641: coeff = 24'd13532841;
            12'd2642: coeff = 24'd13522668;
            12'd2643: coeff = 24'd13512483;
            12'd2644: coeff = 24'd13502286;
            12'd2645: coeff = 24'd13492077;
            12'd2646: coeff = 24'd13481856;
            12'd2647: coeff = 24'd13471623;
            12'd2648: coeff = 24'd13461378;
            12'd2649: coeff = 24'd13451121;
            12'd2650: coeff = 24'd13440852;
            12'd2651: coeff = 24'd13430571;
            12'd2652: coeff = 24'd13420278;
            12'd2653: coeff = 24'd13409974;
            12'd2654: coeff = 24'd13399657;
            12'd2655: coeff = 24'd13389329;
            12'd2656: coeff = 24'd13378989;
            12'd2657: coeff = 24'd13368638;
            12'd2658: coeff = 24'd13358274;
            12'd2659: coeff = 24'd13347899;
            12'd2660: coeff = 24'd13337512;
            12'd2661: coeff = 24'd13327114;
            12'd2662: coeff = 24'd13316704;
            12'd2663: coeff = 24'd13306282;
            12'd2664: coeff = 24'd13295849;
            12'd2665: coeff = 24'd13285404;
            12'd2666: coeff = 24'd13274948;
            12'd2667: coeff = 24'd13264480;
            12'd2668: coeff = 24'd13254001;
            12'd2669: coeff = 24'd13243510;
            12'd2670: coeff = 24'd13233008;
            12'd2671: coeff = 24'd13222494;
            12'd2672: coeff = 24'd13211970;
            12'd2673: coeff = 24'd13201433;
            12'd2674: coeff = 24'd13190886;
            12'd2675: coeff = 24'd13180327;
            12'd2676: coeff = 24'd13169756;
            12'd2677: coeff = 24'd13159175;
            12'd2678: coeff = 24'd13148582;
            12'd2679: coeff = 24'd13137978;
            12'd2680: coeff = 24'd13127363;
            12'd2681: coeff = 24'd13116737;
            12'd2682: coeff = 24'd13106100;
            12'd2683: coeff = 24'd13095451;
            12'd2684: coeff = 24'd13084791;
            12'd2685: coeff = 24'd13074121;
            12'd2686: coeff = 24'd13063439;
            12'd2687: coeff = 24'd13052747;
            12'd2688: coeff = 24'd13042043;
            12'd2689: coeff = 24'd13031328;
            12'd2690: coeff = 24'd13020603;
            12'd2691: coeff = 24'd13009866;
            12'd2692: coeff = 24'd12999119;
            12'd2693: coeff = 24'd12988361;
            12'd2694: coeff = 24'd12977592;
            12'd2695: coeff = 24'd12966812;
            12'd2696: coeff = 24'd12956021;
            12'd2697: coeff = 24'd12945220;
            12'd2698: coeff = 24'd12934408;
            12'd2699: coeff = 24'd12923585;
            12'd2700: coeff = 24'd12912752;
            12'd2701: coeff = 24'd12901908;
            12'd2702: coeff = 24'd12891053;
            12'd2703: coeff = 24'd12880188;
            12'd2704: coeff = 24'd12869312;
            12'd2705: coeff = 24'd12858425;
            12'd2706: coeff = 24'd12847528;
            12'd2707: coeff = 24'd12836621;
            12'd2708: coeff = 24'd12825703;
            12'd2709: coeff = 24'd12814775;
            12'd2710: coeff = 24'd12803836;
            12'd2711: coeff = 24'd12792887;
            12'd2712: coeff = 24'd12781927;
            12'd2713: coeff = 24'd12770957;
            12'd2714: coeff = 24'd12759977;
            12'd2715: coeff = 24'd12748986;
            12'd2716: coeff = 24'd12737986;
            12'd2717: coeff = 24'd12726975;
            12'd2718: coeff = 24'd12715953;
            12'd2719: coeff = 24'd12704922;
            12'd2720: coeff = 24'd12693880;
            12'd2721: coeff = 24'd12682829;
            12'd2722: coeff = 24'd12671767;
            12'd2723: coeff = 24'd12660695;
            12'd2724: coeff = 24'd12649613;
            12'd2725: coeff = 24'd12638521;
            12'd2726: coeff = 24'd12627419;
            12'd2727: coeff = 24'd12616307;
            12'd2728: coeff = 24'd12605185;
            12'd2729: coeff = 24'd12594053;
            12'd2730: coeff = 24'd12582912;
            12'd2731: coeff = 24'd12571760;
            12'd2732: coeff = 24'd12560598;
            12'd2733: coeff = 24'd12549427;
            12'd2734: coeff = 24'd12538246;
            12'd2735: coeff = 24'd12527055;
            12'd2736: coeff = 24'd12515854;
            12'd2737: coeff = 24'd12504644;
            12'd2738: coeff = 24'd12493424;
            12'd2739: coeff = 24'd12482194;
            12'd2740: coeff = 24'd12470955;
            12'd2741: coeff = 24'd12459706;
            12'd2742: coeff = 24'd12448448;
            12'd2743: coeff = 24'd12437180;
            12'd2744: coeff = 24'd12425902;
            12'd2745: coeff = 24'd12414615;
            12'd2746: coeff = 24'd12403318;
            12'd2747: coeff = 24'd12392012;
            12'd2748: coeff = 24'd12380697;
            12'd2749: coeff = 24'd12369372;
            12'd2750: coeff = 24'd12358038;
            12'd2751: coeff = 24'd12346694;
            12'd2752: coeff = 24'd12335341;
            12'd2753: coeff = 24'd12323979;
            12'd2754: coeff = 24'd12312608;
            12'd2755: coeff = 24'd12301227;
            12'd2756: coeff = 24'd12289837;
            12'd2757: coeff = 24'd12278438;
            12'd2758: coeff = 24'd12267030;
            12'd2759: coeff = 24'd12255612;
            12'd2760: coeff = 24'd12244186;
            12'd2761: coeff = 24'd12232750;
            12'd2762: coeff = 24'd12221306;
            12'd2763: coeff = 24'd12209852;
            12'd2764: coeff = 24'd12198389;
            12'd2765: coeff = 24'd12186918;
            12'd2766: coeff = 24'd12175437;
            12'd2767: coeff = 24'd12163948;
            12'd2768: coeff = 24'd12152449;
            12'd2769: coeff = 24'd12140942;
            12'd2770: coeff = 24'd12129426;
            12'd2771: coeff = 24'd12117901;
            12'd2772: coeff = 24'd12106368;
            12'd2773: coeff = 24'd12094825;
            12'd2774: coeff = 24'd12083274;
            12'd2775: coeff = 24'd12071714;
            12'd2776: coeff = 24'd12060146;
            12'd2777: coeff = 24'd12048569;
            12'd2778: coeff = 24'd12036983;
            12'd2779: coeff = 24'd12025389;
            12'd2780: coeff = 24'd12013786;
            12'd2781: coeff = 24'd12002174;
            12'd2782: coeff = 24'd11990554;
            12'd2783: coeff = 24'd11978926;
            12'd2784: coeff = 24'd11967289;
            12'd2785: coeff = 24'd11955644;
            12'd2786: coeff = 24'd11943990;
            12'd2787: coeff = 24'd11932328;
            12'd2788: coeff = 24'd11920658;
            12'd2789: coeff = 24'd11908979;
            12'd2790: coeff = 24'd11897292;
            12'd2791: coeff = 24'd11885597;
            12'd2792: coeff = 24'd11873893;
            12'd2793: coeff = 24'd11862182;
            12'd2794: coeff = 24'd11850462;
            12'd2795: coeff = 24'd11838734;
            12'd2796: coeff = 24'd11826998;
            12'd2797: coeff = 24'd11815253;
            12'd2798: coeff = 24'd11803501;
            12'd2799: coeff = 24'd11791741;
            12'd2800: coeff = 24'd11779972;
            12'd2801: coeff = 24'd11768196;
            12'd2802: coeff = 24'd11756412;
            12'd2803: coeff = 24'd11744620;
            12'd2804: coeff = 24'd11732819;
            12'd2805: coeff = 24'd11721011;
            12'd2806: coeff = 24'd11709196;
            12'd2807: coeff = 24'd11697372;
            12'd2808: coeff = 24'd11685540;
            12'd2809: coeff = 24'd11673701;
            12'd2810: coeff = 24'd11661854;
            12'd2811: coeff = 24'd11650000;
            12'd2812: coeff = 24'd11638137;
            12'd2813: coeff = 24'd11626267;
            12'd2814: coeff = 24'd11614390;
            12'd2815: coeff = 24'd11602504;
            12'd2816: coeff = 24'd11590612;
            12'd2817: coeff = 24'd11578711;
            12'd2818: coeff = 24'd11566804;
            12'd2819: coeff = 24'd11554888;
            12'd2820: coeff = 24'd11542966;
            12'd2821: coeff = 24'd11531035;
            12'd2822: coeff = 24'd11519098;
            12'd2823: coeff = 24'd11507153;
            12'd2824: coeff = 24'd11495201;
            12'd2825: coeff = 24'd11483241;
            12'd2826: coeff = 24'd11471274;
            12'd2827: coeff = 24'd11459300;
            12'd2828: coeff = 24'd11447319;
            12'd2829: coeff = 24'd11435330;
            12'd2830: coeff = 24'd11423334;
            12'd2831: coeff = 24'd11411331;
            12'd2832: coeff = 24'd11399321;
            12'd2833: coeff = 24'd11387304;
            12'd2834: coeff = 24'd11375280;
            12'd2835: coeff = 24'd11363249;
            12'd2836: coeff = 24'd11351211;
            12'd2837: coeff = 24'd11339166;
            12'd2838: coeff = 24'd11327113;
            12'd2839: coeff = 24'd11315054;
            12'd2840: coeff = 24'd11302988;
            12'd2841: coeff = 24'd11290916;
            12'd2842: coeff = 24'd11278836;
            12'd2843: coeff = 24'd11266750;
            12'd2844: coeff = 24'd11254656;
            12'd2845: coeff = 24'd11242557;
            12'd2846: coeff = 24'd11230450;
            12'd2847: coeff = 24'd11218337;
            12'd2848: coeff = 24'd11206217;
            12'd2849: coeff = 24'd11194090;
            12'd2850: coeff = 24'd11181957;
            12'd2851: coeff = 24'd11169817;
            12'd2852: coeff = 24'd11157670;
            12'd2853: coeff = 24'd11145518;
            12'd2854: coeff = 24'd11133358;
            12'd2855: coeff = 24'd11121192;
            12'd2856: coeff = 24'd11109020;
            12'd2857: coeff = 24'd11096841;
            12'd2858: coeff = 24'd11084656;
            12'd2859: coeff = 24'd11072465;
            12'd2860: coeff = 24'd11060267;
            12'd2861: coeff = 24'd11048063;
            12'd2862: coeff = 24'd11035853;
            12'd2863: coeff = 24'd11023636;
            12'd2864: coeff = 24'd11011414;
            12'd2865: coeff = 24'd10999185;
            12'd2866: coeff = 24'd10986950;
            12'd2867: coeff = 24'd10974709;
            12'd2868: coeff = 24'd10962461;
            12'd2869: coeff = 24'd10950208;
            12'd2870: coeff = 24'd10937949;
            12'd2871: coeff = 24'd10925683;
            12'd2872: coeff = 24'd10913412;
            12'd2873: coeff = 24'd10901135;
            12'd2874: coeff = 24'd10888852;
            12'd2875: coeff = 24'd10876563;
            12'd2876: coeff = 24'd10864268;
            12'd2877: coeff = 24'd10851967;
            12'd2878: coeff = 24'd10839660;
            12'd2879: coeff = 24'd10827348;
            12'd2880: coeff = 24'd10815030;
            12'd2881: coeff = 24'd10802706;
            12'd2882: coeff = 24'd10790377;
            12'd2883: coeff = 24'd10778042;
            12'd2884: coeff = 24'd10765701;
            12'd2885: coeff = 24'd10753355;
            12'd2886: coeff = 24'd10741003;
            12'd2887: coeff = 24'd10728646;
            12'd2888: coeff = 24'd10716283;
            12'd2889: coeff = 24'd10703914;
            12'd2890: coeff = 24'd10691540;
            12'd2891: coeff = 24'd10679161;
            12'd2892: coeff = 24'd10666776;
            12'd2893: coeff = 24'd10654386;
            12'd2894: coeff = 24'd10641991;
            12'd2895: coeff = 24'd10629590;
            12'd2896: coeff = 24'd10617184;
            12'd2897: coeff = 24'd10604773;
            12'd2898: coeff = 24'd10592357;
            12'd2899: coeff = 24'd10579935;
            12'd2900: coeff = 24'd10567508;
            12'd2901: coeff = 24'd10555076;
            12'd2902: coeff = 24'd10542639;
            12'd2903: coeff = 24'd10530197;
            12'd2904: coeff = 24'd10517750;
            12'd2905: coeff = 24'd10505298;
            12'd2906: coeff = 24'd10492841;
            12'd2907: coeff = 24'd10480379;
            12'd2908: coeff = 24'd10467912;
            12'd2909: coeff = 24'd10455440;
            12'd2910: coeff = 24'd10442963;
            12'd2911: coeff = 24'd10430482;
            12'd2912: coeff = 24'd10417995;
            12'd2913: coeff = 24'd10405504;
            12'd2914: coeff = 24'd10393008;
            12'd2915: coeff = 24'd10380508;
            12'd2916: coeff = 24'd10368002;
            12'd2917: coeff = 24'd10355492;
            12'd2918: coeff = 24'd10342978;
            12'd2919: coeff = 24'd10330459;
            12'd2920: coeff = 24'd10317935;
            12'd2921: coeff = 24'd10305407;
            12'd2922: coeff = 24'd10292874;
            12'd2923: coeff = 24'd10280336;
            12'd2924: coeff = 24'd10267795;
            12'd2925: coeff = 24'd10255248;
            12'd2926: coeff = 24'd10242698;
            12'd2927: coeff = 24'd10230143;
            12'd2928: coeff = 24'd10217584;
            12'd2929: coeff = 24'd10205020;
            12'd2930: coeff = 24'd10192452;
            12'd2931: coeff = 24'd10179880;
            12'd2932: coeff = 24'd10167304;
            12'd2933: coeff = 24'd10154723;
            12'd2934: coeff = 24'd10142138;
            12'd2935: coeff = 24'd10129550;
            12'd2936: coeff = 24'd10116957;
            12'd2937: coeff = 24'd10104360;
            12'd2938: coeff = 24'd10091759;
            12'd2939: coeff = 24'd10079154;
            12'd2940: coeff = 24'd10066545;
            12'd2941: coeff = 24'd10053932;
            12'd2942: coeff = 24'd10041315;
            12'd2943: coeff = 24'd10028694;
            12'd2944: coeff = 24'd10016069;
            12'd2945: coeff = 24'd10003441;
            12'd2946: coeff = 24'd9990809;
            12'd2947: coeff = 24'd9978173;
            12'd2948: coeff = 24'd9965533;
            12'd2949: coeff = 24'd9952889;
            12'd2950: coeff = 24'd9940242;
            12'd2951: coeff = 24'd9927591;
            12'd2952: coeff = 24'd9914937;
            12'd2953: coeff = 24'd9902279;
            12'd2954: coeff = 24'd9889617;
            12'd2955: coeff = 24'd9876952;
            12'd2956: coeff = 24'd9864283;
            12'd2957: coeff = 24'd9851611;
            12'd2958: coeff = 24'd9838936;
            12'd2959: coeff = 24'd9826257;
            12'd2960: coeff = 24'd9813574;
            12'd2961: coeff = 24'd9800889;
            12'd2962: coeff = 24'd9788200;
            12'd2963: coeff = 24'd9775507;
            12'd2964: coeff = 24'd9762812;
            12'd2965: coeff = 24'd9750113;
            12'd2966: coeff = 24'd9737411;
            12'd2967: coeff = 24'd9724706;
            12'd2968: coeff = 24'd9711997;
            12'd2969: coeff = 24'd9699286;
            12'd2970: coeff = 24'd9686571;
            12'd2971: coeff = 24'd9673854;
            12'd2972: coeff = 24'd9661133;
            12'd2973: coeff = 24'd9648409;
            12'd2974: coeff = 24'd9635683;
            12'd2975: coeff = 24'd9622953;
            12'd2976: coeff = 24'd9610221;
            12'd2977: coeff = 24'd9597485;
            12'd2978: coeff = 24'd9584747;
            12'd2979: coeff = 24'd9572006;
            12'd2980: coeff = 24'd9559262;
            12'd2981: coeff = 24'd9546516;
            12'd2982: coeff = 24'd9533767;
            12'd2983: coeff = 24'd9521015;
            12'd2984: coeff = 24'd9508260;
            12'd2985: coeff = 24'd9495503;
            12'd2986: coeff = 24'd9482743;
            12'd2987: coeff = 24'd9469981;
            12'd2988: coeff = 24'd9457216;
            12'd2989: coeff = 24'd9444448;
            12'd2990: coeff = 24'd9431678;
            12'd2991: coeff = 24'd9418906;
            12'd2992: coeff = 24'd9406131;
            12'd2993: coeff = 24'd9393354;
            12'd2994: coeff = 24'd9380574;
            12'd2995: coeff = 24'd9367792;
            12'd2996: coeff = 24'd9355008;
            12'd2997: coeff = 24'd9342221;
            12'd2998: coeff = 24'd9329432;
            12'd2999: coeff = 24'd9316641;
            12'd3000: coeff = 24'd9303848;
            12'd3001: coeff = 24'd9291053;
            12'd3002: coeff = 24'd9278255;
            12'd3003: coeff = 24'd9265456;
            12'd3004: coeff = 24'd9252654;
            12'd3005: coeff = 24'd9239851;
            12'd3006: coeff = 24'd9227045;
            12'd3007: coeff = 24'd9214237;
            12'd3008: coeff = 24'd9201428;
            12'd3009: coeff = 24'd9188616;
            12'd3010: coeff = 24'd9175803;
            12'd3011: coeff = 24'd9162988;
            12'd3012: coeff = 24'd9150170;
            12'd3013: coeff = 24'd9137352;
            12'd3014: coeff = 24'd9124531;
            12'd3015: coeff = 24'd9111709;
            12'd3016: coeff = 24'd9098885;
            12'd3017: coeff = 24'd9086059;
            12'd3018: coeff = 24'd9073232;
            12'd3019: coeff = 24'd9060403;
            12'd3020: coeff = 24'd9047572;
            12'd3021: coeff = 24'd9034740;
            12'd3022: coeff = 24'd9021906;
            12'd3023: coeff = 24'd9009071;
            12'd3024: coeff = 24'd8996235;
            12'd3025: coeff = 24'd8983397;
            12'd3026: coeff = 24'd8970557;
            12'd3027: coeff = 24'd8957716;
            12'd3028: coeff = 24'd8944874;
            12'd3029: coeff = 24'd8932031;
            12'd3030: coeff = 24'd8919186;
            12'd3031: coeff = 24'd8906340;
            12'd3032: coeff = 24'd8893493;
            12'd3033: coeff = 24'd8880645;
            12'd3034: coeff = 24'd8867795;
            12'd3035: coeff = 24'd8854945;
            12'd3036: coeff = 24'd8842093;
            12'd3037: coeff = 24'd8829240;
            12'd3038: coeff = 24'd8816386;
            12'd3039: coeff = 24'd8803531;
            12'd3040: coeff = 24'd8790675;
            12'd3041: coeff = 24'd8777819;
            12'd3042: coeff = 24'd8764961;
            12'd3043: coeff = 24'd8752102;
            12'd3044: coeff = 24'd8739243;
            12'd3045: coeff = 24'd8726383;
            12'd3046: coeff = 24'd8713522;
            12'd3047: coeff = 24'd8700660;
            12'd3048: coeff = 24'd8687797;
            12'd3049: coeff = 24'd8674934;
            12'd3050: coeff = 24'd8662070;
            12'd3051: coeff = 24'd8649205;
            12'd3052: coeff = 24'd8636340;
            12'd3053: coeff = 24'd8623474;
            12'd3054: coeff = 24'd8610608;
            12'd3055: coeff = 24'd8597741;
            12'd3056: coeff = 24'd8584874;
            12'd3057: coeff = 24'd8572006;
            12'd3058: coeff = 24'd8559138;
            12'd3059: coeff = 24'd8546269;
            12'd3060: coeff = 24'd8533400;
            12'd3061: coeff = 24'd8520531;
            12'd3062: coeff = 24'd8507661;
            12'd3063: coeff = 24'd8494791;
            12'd3064: coeff = 24'd8481921;
            12'd3065: coeff = 24'd8469051;
            12'd3066: coeff = 24'd8456180;
            12'd3067: coeff = 24'd8443309;
            12'd3068: coeff = 24'd8430438;
            12'd3069: coeff = 24'd8417567;
            12'd3070: coeff = 24'd8404696;
            12'd3071: coeff = 24'd8391825;
            12'd3072: coeff = 24'd8378954;
            12'd3073: coeff = 24'd8366083;
            12'd3074: coeff = 24'd8353212;
            12'd3075: coeff = 24'd8340341;
            12'd3076: coeff = 24'd8327470;
            12'd3077: coeff = 24'd8314600;
            12'd3078: coeff = 24'd8301729;
            12'd3079: coeff = 24'd8288859;
            12'd3080: coeff = 24'd8275989;
            12'd3081: coeff = 24'd8263119;
            12'd3082: coeff = 24'd8250249;
            12'd3083: coeff = 24'd8237380;
            12'd3084: coeff = 24'd8224511;
            12'd3085: coeff = 24'd8211643;
            12'd3086: coeff = 24'd8198775;
            12'd3087: coeff = 24'd8185907;
            12'd3088: coeff = 24'd8173040;
            12'd3089: coeff = 24'd8160174;
            12'd3090: coeff = 24'd8147308;
            12'd3091: coeff = 24'd8134442;
            12'd3092: coeff = 24'd8121577;
            12'd3093: coeff = 24'd8108713;
            12'd3094: coeff = 24'd8095849;
            12'd3095: coeff = 24'd8082986;
            12'd3096: coeff = 24'd8070124;
            12'd3097: coeff = 24'd8057263;
            12'd3098: coeff = 24'd8044402;
            12'd3099: coeff = 24'd8031542;
            12'd3100: coeff = 24'd8018683;
            12'd3101: coeff = 24'd8005825;
            12'd3102: coeff = 24'd7992968;
            12'd3103: coeff = 24'd7980112;
            12'd3104: coeff = 24'd7967256;
            12'd3105: coeff = 24'd7954402;
            12'd3106: coeff = 24'd7941548;
            12'd3107: coeff = 24'd7928696;
            12'd3108: coeff = 24'd7915845;
            12'd3109: coeff = 24'd7902995;
            12'd3110: coeff = 24'd7890146;
            12'd3111: coeff = 24'd7877298;
            12'd3112: coeff = 24'd7864452;
            12'd3113: coeff = 24'd7851606;
            12'd3114: coeff = 24'd7838762;
            12'd3115: coeff = 24'd7825919;
            12'd3116: coeff = 24'd7813078;
            12'd3117: coeff = 24'd7800238;
            12'd3118: coeff = 24'd7787399;
            12'd3119: coeff = 24'd7774562;
            12'd3120: coeff = 24'd7761726;
            12'd3121: coeff = 24'd7748892;
            12'd3122: coeff = 24'd7736059;
            12'd3123: coeff = 24'd7723227;
            12'd3124: coeff = 24'd7710398;
            12'd3125: coeff = 24'd7697570;
            12'd3126: coeff = 24'd7684743;
            12'd3127: coeff = 24'd7671918;
            12'd3128: coeff = 24'd7659095;
            12'd3129: coeff = 24'd7646273;
            12'd3130: coeff = 24'd7633454;
            12'd3131: coeff = 24'd7620636;
            12'd3132: coeff = 24'd7607820;
            12'd3133: coeff = 24'd7595005;
            12'd3134: coeff = 24'd7582193;
            12'd3135: coeff = 24'd7569382;
            12'd3136: coeff = 24'd7556574;
            12'd3137: coeff = 24'd7543767;
            12'd3138: coeff = 24'd7530962;
            12'd3139: coeff = 24'd7518160;
            12'd3140: coeff = 24'd7505359;
            12'd3141: coeff = 24'd7492561;
            12'd3142: coeff = 24'd7479764;
            12'd3143: coeff = 24'd7466970;
            12'd3144: coeff = 24'd7454178;
            12'd3145: coeff = 24'd7441388;
            12'd3146: coeff = 24'd7428600;
            12'd3147: coeff = 24'd7415815;
            12'd3148: coeff = 24'd7403032;
            12'd3149: coeff = 24'd7390251;
            12'd3150: coeff = 24'd7377473;
            12'd3151: coeff = 24'd7364696;
            12'd3152: coeff = 24'd7351923;
            12'd3153: coeff = 24'd7339152;
            12'd3154: coeff = 24'd7326383;
            12'd3155: coeff = 24'd7313617;
            12'd3156: coeff = 24'd7300853;
            12'd3157: coeff = 24'd7288092;
            12'd3158: coeff = 24'd7275333;
            12'd3159: coeff = 24'd7262577;
            12'd3160: coeff = 24'd7249824;
            12'd3161: coeff = 24'd7237073;
            12'd3162: coeff = 24'd7224325;
            12'd3163: coeff = 24'd7211580;
            12'd3164: coeff = 24'd7198838;
            12'd3165: coeff = 24'd7186098;
            12'd3166: coeff = 24'd7173362;
            12'd3167: coeff = 24'd7160628;
            12'd3168: coeff = 24'd7147897;
            12'd3169: coeff = 24'd7135169;
            12'd3170: coeff = 24'd7122443;
            12'd3171: coeff = 24'd7109721;
            12'd3172: coeff = 24'd7097002;
            12'd3173: coeff = 24'd7084286;
            12'd3174: coeff = 24'd7071573;
            12'd3175: coeff = 24'd7058863;
            12'd3176: coeff = 24'd7046156;
            12'd3177: coeff = 24'd7033453;
            12'd3178: coeff = 24'd7020752;
            12'd3179: coeff = 24'd7008055;
            12'd3180: coeff = 24'd6995361;
            12'd3181: coeff = 24'd6982670;
            12'd3182: coeff = 24'd6969983;
            12'd3183: coeff = 24'd6957299;
            12'd3184: coeff = 24'd6944618;
            12'd3185: coeff = 24'd6931941;
            12'd3186: coeff = 24'd6919267;
            12'd3187: coeff = 24'd6906597;
            12'd3188: coeff = 24'd6893930;
            12'd3189: coeff = 24'd6881267;
            12'd3190: coeff = 24'd6868607;
            12'd3191: coeff = 24'd6855950;
            12'd3192: coeff = 24'd6843298;
            12'd3193: coeff = 24'd6830649;
            12'd3194: coeff = 24'd6818003;
            12'd3195: coeff = 24'd6805362;
            12'd3196: coeff = 24'd6792724;
            12'd3197: coeff = 24'd6780090;
            12'd3198: coeff = 24'd6767459;
            12'd3199: coeff = 24'd6754833;
            12'd3200: coeff = 24'd6742210;
            12'd3201: coeff = 24'd6729591;
            12'd3202: coeff = 24'd6716976;
            12'd3203: coeff = 24'd6704365;
            12'd3204: coeff = 24'd6691758;
            12'd3205: coeff = 24'd6679155;
            12'd3206: coeff = 24'd6666556;
            12'd3207: coeff = 24'd6653961;
            12'd3208: coeff = 24'd6641370;
            12'd3209: coeff = 24'd6628784;
            12'd3210: coeff = 24'd6616201;
            12'd3211: coeff = 24'd6603623;
            12'd3212: coeff = 24'd6591048;
            12'd3213: coeff = 24'd6578478;
            12'd3214: coeff = 24'd6565913;
            12'd3215: coeff = 24'd6553351;
            12'd3216: coeff = 24'd6540794;
            12'd3217: coeff = 24'd6528241;
            12'd3218: coeff = 24'd6515693;
            12'd3219: coeff = 24'd6503149;
            12'd3220: coeff = 24'd6490609;
            12'd3221: coeff = 24'd6478074;
            12'd3222: coeff = 24'd6465544;
            12'd3223: coeff = 24'd6453018;
            12'd3224: coeff = 24'd6440496;
            12'd3225: coeff = 24'd6427979;
            12'd3226: coeff = 24'd6415467;
            12'd3227: coeff = 24'd6402959;
            12'd3228: coeff = 24'd6390456;
            12'd3229: coeff = 24'd6377958;
            12'd3230: coeff = 24'd6365465;
            12'd3231: coeff = 24'd6352976;
            12'd3232: coeff = 24'd6340492;
            12'd3233: coeff = 24'd6328013;
            12'd3234: coeff = 24'd6315538;
            12'd3235: coeff = 24'd6303069;
            12'd3236: coeff = 24'd6290604;
            12'd3237: coeff = 24'd6278145;
            12'd3238: coeff = 24'd6265690;
            12'd3239: coeff = 24'd6253241;
            12'd3240: coeff = 24'd6240796;
            12'd3241: coeff = 24'd6228356;
            12'd3242: coeff = 24'd6215922;
            12'd3243: coeff = 24'd6203493;
            12'd3244: coeff = 24'd6191068;
            12'd3245: coeff = 24'd6178649;
            12'd3246: coeff = 24'd6166236;
            12'd3247: coeff = 24'd6153827;
            12'd3248: coeff = 24'd6141424;
            12'd3249: coeff = 24'd6129026;
            12'd3250: coeff = 24'd6116633;
            12'd3251: coeff = 24'd6104246;
            12'd3252: coeff = 24'd6091864;
            12'd3253: coeff = 24'd6079487;
            12'd3254: coeff = 24'd6067116;
            12'd3255: coeff = 24'd6054750;
            12'd3256: coeff = 24'd6042390;
            12'd3257: coeff = 24'd6030035;
            12'd3258: coeff = 24'd6017686;
            12'd3259: coeff = 24'd6005343;
            12'd3260: coeff = 24'd5993005;
            12'd3261: coeff = 24'd5980673;
            12'd3262: coeff = 24'd5968346;
            12'd3263: coeff = 24'd5956025;
            12'd3264: coeff = 24'd5943710;
            12'd3265: coeff = 24'd5931401;
            12'd3266: coeff = 24'd5919097;
            12'd3267: coeff = 24'd5906799;
            12'd3268: coeff = 24'd5894507;
            12'd3269: coeff = 24'd5882221;
            12'd3270: coeff = 24'd5869941;
            12'd3271: coeff = 24'd5857666;
            12'd3272: coeff = 24'd5845398;
            12'd3273: coeff = 24'd5833136;
            12'd3274: coeff = 24'd5820880;
            12'd3275: coeff = 24'd5808629;
            12'd3276: coeff = 24'd5796385;
            12'd3277: coeff = 24'd5784147;
            12'd3278: coeff = 24'd5771915;
            12'd3279: coeff = 24'd5759689;
            12'd3280: coeff = 24'd5747470;
            12'd3281: coeff = 24'd5735256;
            12'd3282: coeff = 24'd5723049;
            12'd3283: coeff = 24'd5710848;
            12'd3284: coeff = 24'd5698654;
            12'd3285: coeff = 24'd5686465;
            12'd3286: coeff = 24'd5674284;
            12'd3287: coeff = 24'd5662108;
            12'd3288: coeff = 24'd5649939;
            12'd3289: coeff = 24'd5637776;
            12'd3290: coeff = 24'd5625620;
            12'd3291: coeff = 24'd5613471;
            12'd3292: coeff = 24'd5601327;
            12'd3293: coeff = 24'd5589191;
            12'd3294: coeff = 24'd5577061;
            12'd3295: coeff = 24'd5564938;
            12'd3296: coeff = 24'd5552821;
            12'd3297: coeff = 24'd5540711;
            12'd3298: coeff = 24'd5528608;
            12'd3299: coeff = 24'd5516511;
            12'd3300: coeff = 24'd5504421;
            12'd3301: coeff = 24'd5492338;
            12'd3302: coeff = 24'd5480262;
            12'd3303: coeff = 24'd5468193;
            12'd3304: coeff = 24'd5456130;
            12'd3305: coeff = 24'd5444075;
            12'd3306: coeff = 24'd5432026;
            12'd3307: coeff = 24'd5419984;
            12'd3308: coeff = 24'd5407950;
            12'd3309: coeff = 24'd5395922;
            12'd3310: coeff = 24'd5383901;
            12'd3311: coeff = 24'd5371888;
            12'd3312: coeff = 24'd5359881;
            12'd3313: coeff = 24'd5347882;
            12'd3314: coeff = 24'd5335890;
            12'd3315: coeff = 24'd5323905;
            12'd3316: coeff = 24'd5311927;
            12'd3317: coeff = 24'd5299957;
            12'd3318: coeff = 24'd5287993;
            12'd3319: coeff = 24'd5276037;
            12'd3320: coeff = 24'd5264089;
            12'd3321: coeff = 24'd5252147;
            12'd3322: coeff = 24'd5240214;
            12'd3323: coeff = 24'd5228287;
            12'd3324: coeff = 24'd5216368;
            12'd3325: coeff = 24'd5204457;
            12'd3326: coeff = 24'd5192552;
            12'd3327: coeff = 24'd5180656;
            12'd3328: coeff = 24'd5168767;
            12'd3329: coeff = 24'd5156886;
            12'd3330: coeff = 24'd5145012;
            12'd3331: coeff = 24'd5133146;
            12'd3332: coeff = 24'd5121287;
            12'd3333: coeff = 24'd5109436;
            12'd3334: coeff = 24'd5097593;
            12'd3335: coeff = 24'd5085758;
            12'd3336: coeff = 24'd5073930;
            12'd3337: coeff = 24'd5062111;
            12'd3338: coeff = 24'd5050299;
            12'd3339: coeff = 24'd5038495;
            12'd3340: coeff = 24'd5026698;
            12'd3341: coeff = 24'd5014910;
            12'd3342: coeff = 24'd5003130;
            12'd3343: coeff = 24'd4991357;
            12'd3344: coeff = 24'd4979593;
            12'd3345: coeff = 24'd4967837;
            12'd3346: coeff = 24'd4956088;
            12'd3347: coeff = 24'd4944348;
            12'd3348: coeff = 24'd4932616;
            12'd3349: coeff = 24'd4920892;
            12'd3350: coeff = 24'd4909176;
            12'd3351: coeff = 24'd4897469;
            12'd3352: coeff = 24'd4885769;
            12'd3353: coeff = 24'd4874078;
            12'd3354: coeff = 24'd4862395;
            12'd3355: coeff = 24'd4850721;
            12'd3356: coeff = 24'd4839055;
            12'd3357: coeff = 24'd4827397;
            12'd3358: coeff = 24'd4815747;
            12'd3359: coeff = 24'd4804106;
            12'd3360: coeff = 24'd4792474;
            12'd3361: coeff = 24'd4780849;
            12'd3362: coeff = 24'd4769234;
            12'd3363: coeff = 24'd4757627;
            12'd3364: coeff = 24'd4746028;
            12'd3365: coeff = 24'd4734438;
            12'd3366: coeff = 24'd4722857;
            12'd3367: coeff = 24'd4711284;
            12'd3368: coeff = 24'd4699720;
            12'd3369: coeff = 24'd4688164;
            12'd3370: coeff = 24'd4676617;
            12'd3371: coeff = 24'd4665079;
            12'd3372: coeff = 24'd4653550;
            12'd3373: coeff = 24'd4642030;
            12'd3374: coeff = 24'd4630518;
            12'd3375: coeff = 24'd4619015;
            12'd3376: coeff = 24'd4607521;
            12'd3377: coeff = 24'd4596036;
            12'd3378: coeff = 24'd4584560;
            12'd3379: coeff = 24'd4573093;
            12'd3380: coeff = 24'd4561635;
            12'd3381: coeff = 24'd4550186;
            12'd3382: coeff = 24'd4538746;
            12'd3383: coeff = 24'd4527315;
            12'd3384: coeff = 24'd4515893;
            12'd3385: coeff = 24'd4504480;
            12'd3386: coeff = 24'd4493076;
            12'd3387: coeff = 24'd4481682;
            12'd3388: coeff = 24'd4470297;
            12'd3389: coeff = 24'd4458921;
            12'd3390: coeff = 24'd4447554;
            12'd3391: coeff = 24'd4436196;
            12'd3392: coeff = 24'd4424848;
            12'd3393: coeff = 24'd4413509;
            12'd3394: coeff = 24'd4402179;
            12'd3395: coeff = 24'd4390859;
            12'd3396: coeff = 24'd4379549;
            12'd3397: coeff = 24'd4368247;
            12'd3398: coeff = 24'd4356955;
            12'd3399: coeff = 24'd4345673;
            12'd3400: coeff = 24'd4334400;
            12'd3401: coeff = 24'd4323137;
            12'd3402: coeff = 24'd4311883;
            12'd3403: coeff = 24'd4300639;
            12'd3404: coeff = 24'd4289405;
            12'd3405: coeff = 24'd4278180;
            12'd3406: coeff = 24'd4266964;
            12'd3407: coeff = 24'd4255759;
            12'd3408: coeff = 24'd4244563;
            12'd3409: coeff = 24'd4233377;
            12'd3410: coeff = 24'd4222201;
            12'd3411: coeff = 24'd4211035;
            12'd3412: coeff = 24'd4199878;
            12'd3413: coeff = 24'd4188731;
            12'd3414: coeff = 24'd4177595;
            12'd3415: coeff = 24'd4166468;
            12'd3416: coeff = 24'd4155351;
            12'd3417: coeff = 24'd4144244;
            12'd3418: coeff = 24'd4133147;
            12'd3419: coeff = 24'd4122060;
            12'd3420: coeff = 24'd4110983;
            12'd3421: coeff = 24'd4099916;
            12'd3422: coeff = 24'd4088859;
            12'd3423: coeff = 24'd4077812;
            12'd3424: coeff = 24'd4066776;
            12'd3425: coeff = 24'd4055750;
            12'd3426: coeff = 24'd4044734;
            12'd3427: coeff = 24'd4033728;
            12'd3428: coeff = 24'd4022732;
            12'd3429: coeff = 24'd4011747;
            12'd3430: coeff = 24'd4000772;
            12'd3431: coeff = 24'd3989807;
            12'd3432: coeff = 24'd3978852;
            12'd3433: coeff = 24'd3967908;
            12'd3434: coeff = 24'd3956975;
            12'd3435: coeff = 24'd3946052;
            12'd3436: coeff = 24'd3935139;
            12'd3437: coeff = 24'd3924237;
            12'd3438: coeff = 24'd3913345;
            12'd3439: coeff = 24'd3902464;
            12'd3440: coeff = 24'd3891593;
            12'd3441: coeff = 24'd3880733;
            12'd3442: coeff = 24'd3869884;
            12'd3443: coeff = 24'd3859045;
            12'd3444: coeff = 24'd3848217;
            12'd3445: coeff = 24'd3837400;
            12'd3446: coeff = 24'd3826593;
            12'd3447: coeff = 24'd3815797;
            12'd3448: coeff = 24'd3805012;
            12'd3449: coeff = 24'd3794237;
            12'd3450: coeff = 24'd3783474;
            12'd3451: coeff = 24'd3772721;
            12'd3452: coeff = 24'd3761979;
            12'd3453: coeff = 24'd3751248;
            12'd3454: coeff = 24'd3740528;
            12'd3455: coeff = 24'd3729819;
            12'd3456: coeff = 24'd3719121;
            12'd3457: coeff = 24'd3708434;
            12'd3458: coeff = 24'd3697757;
            12'd3459: coeff = 24'd3687092;
            12'd3460: coeff = 24'd3676438;
            12'd3461: coeff = 24'd3665795;
            12'd3462: coeff = 24'd3655164;
            12'd3463: coeff = 24'd3644543;
            12'd3464: coeff = 24'd3633933;
            12'd3465: coeff = 24'd3623335;
            12'd3466: coeff = 24'd3612748;
            12'd3467: coeff = 24'd3602172;
            12'd3468: coeff = 24'd3591607;
            12'd3469: coeff = 24'd3581054;
            12'd3470: coeff = 24'd3570512;
            12'd3471: coeff = 24'd3559982;
            12'd3472: coeff = 24'd3549462;
            12'd3473: coeff = 24'd3538954;
            12'd3474: coeff = 24'd3528458;
            12'd3475: coeff = 24'd3517973;
            12'd3476: coeff = 24'd3507499;
            12'd3477: coeff = 24'd3497037;
            12'd3478: coeff = 24'd3486587;
            12'd3479: coeff = 24'd3476148;
            12'd3480: coeff = 24'd3465720;
            12'd3481: coeff = 24'd3455305;
            12'd3482: coeff = 24'd3444900;
            12'd3483: coeff = 24'd3434508;
            12'd3484: coeff = 24'd3424127;
            12'd3485: coeff = 24'd3413758;
            12'd3486: coeff = 24'd3403400;
            12'd3487: coeff = 24'd3393054;
            12'd3488: coeff = 24'd3382720;
            12'd3489: coeff = 24'd3372398;
            12'd3490: coeff = 24'd3362088;
            12'd3491: coeff = 24'd3351789;
            12'd3492: coeff = 24'd3341502;
            12'd3493: coeff = 24'd3331227;
            12'd3494: coeff = 24'd3320964;
            12'd3495: coeff = 24'd3310713;
            12'd3496: coeff = 24'd3300474;
            12'd3497: coeff = 24'd3290247;
            12'd3498: coeff = 24'd3280032;
            12'd3499: coeff = 24'd3269829;
            12'd3500: coeff = 24'd3259638;
            12'd3501: coeff = 24'd3249459;
            12'd3502: coeff = 24'd3239292;
            12'd3503: coeff = 24'd3229138;
            12'd3504: coeff = 24'd3218995;
            12'd3505: coeff = 24'd3208865;
            12'd3506: coeff = 24'd3198746;
            12'd3507: coeff = 24'd3188640;
            12'd3508: coeff = 24'd3178547;
            12'd3509: coeff = 24'd3168465;
            12'd3510: coeff = 24'd3158396;
            12'd3511: coeff = 24'd3148339;
            12'd3512: coeff = 24'd3138295;
            12'd3513: coeff = 24'd3128262;
            12'd3514: coeff = 24'd3118243;
            12'd3515: coeff = 24'd3108235;
            12'd3516: coeff = 24'd3098240;
            12'd3517: coeff = 24'd3088258;
            12'd3518: coeff = 24'd3078288;
            12'd3519: coeff = 24'd3068330;
            12'd3520: coeff = 24'd3058385;
            12'd3521: coeff = 24'd3048453;
            12'd3522: coeff = 24'd3038533;
            12'd3523: coeff = 24'd3028626;
            12'd3524: coeff = 24'd3018731;
            12'd3525: coeff = 24'd3008849;
            12'd3526: coeff = 24'd2998980;
            12'd3527: coeff = 24'd2989123;
            12'd3528: coeff = 24'd2979279;
            12'd3529: coeff = 24'd2969448;
            12'd3530: coeff = 24'd2959629;
            12'd3531: coeff = 24'd2949824;
            12'd3532: coeff = 24'd2940031;
            12'd3533: coeff = 24'd2930251;
            12'd3534: coeff = 24'd2920483;
            12'd3535: coeff = 24'd2910729;
            12'd3536: coeff = 24'd2900988;
            12'd3537: coeff = 24'd2891259;
            12'd3538: coeff = 24'd2881544;
            12'd3539: coeff = 24'd2871841;
            12'd3540: coeff = 24'd2862151;
            12'd3541: coeff = 24'd2852475;
            12'd3542: coeff = 24'd2842811;
            12'd3543: coeff = 24'd2833161;
            12'd3544: coeff = 24'd2823523;
            12'd3545: coeff = 24'd2813899;
            12'd3546: coeff = 24'd2804288;
            12'd3547: coeff = 24'd2794690;
            12'd3548: coeff = 24'd2785105;
            12'd3549: coeff = 24'd2775533;
            12'd3550: coeff = 24'd2765975;
            12'd3551: coeff = 24'd2756429;
            12'd3552: coeff = 24'd2746897;
            12'd3553: coeff = 24'd2737379;
            12'd3554: coeff = 24'd2727873;
            12'd3555: coeff = 24'd2718381;
            12'd3556: coeff = 24'd2708903;
            12'd3557: coeff = 24'd2699437;
            12'd3558: coeff = 24'd2689985;
            12'd3559: coeff = 24'd2680547;
            12'd3560: coeff = 24'd2671122;
            12'd3561: coeff = 24'd2661710;
            12'd3562: coeff = 24'd2652312;
            12'd3563: coeff = 24'd2642927;
            12'd3564: coeff = 24'd2633556;
            12'd3565: coeff = 24'd2624198;
            12'd3566: coeff = 24'd2614854;
            12'd3567: coeff = 24'd2605524;
            12'd3568: coeff = 24'd2596207;
            12'd3569: coeff = 24'd2586904;
            12'd3570: coeff = 24'd2577614;
            12'd3571: coeff = 24'd2568339;
            12'd3572: coeff = 24'd2559076;
            12'd3573: coeff = 24'd2549828;
            12'd3574: coeff = 24'd2540593;
            12'd3575: coeff = 24'd2531373;
            12'd3576: coeff = 24'd2522165;
            12'd3577: coeff = 24'd2512972;
            12'd3578: coeff = 24'd2503793;
            12'd3579: coeff = 24'd2494627;
            12'd3580: coeff = 24'd2485475;
            12'd3581: coeff = 24'd2476338;
            12'd3582: coeff = 24'd2467214;
            12'd3583: coeff = 24'd2458104;
            12'd3584: coeff = 24'd2449008;
            12'd3585: coeff = 24'd2439926;
            12'd3586: coeff = 24'd2430858;
            12'd3587: coeff = 24'd2421804;
            12'd3588: coeff = 24'd2412764;
            12'd3589: coeff = 24'd2403738;
            12'd3590: coeff = 24'd2394726;
            12'd3591: coeff = 24'd2385728;
            12'd3592: coeff = 24'd2376745;
            12'd3593: coeff = 24'd2367775;
            12'd3594: coeff = 24'd2358820;
            12'd3595: coeff = 24'd2349879;
            12'd3596: coeff = 24'd2340952;
            12'd3597: coeff = 24'd2332040;
            12'd3598: coeff = 24'd2323141;
            12'd3599: coeff = 24'd2314257;
            12'd3600: coeff = 24'd2305388;
            12'd3601: coeff = 24'd2296532;
            12'd3602: coeff = 24'd2287691;
            12'd3603: coeff = 24'd2278865;
            12'd3604: coeff = 24'd2270052;
            12'd3605: coeff = 24'd2261254;
            12'd3606: coeff = 24'd2252471;
            12'd3607: coeff = 24'd2243702;
            12'd3608: coeff = 24'd2234947;
            12'd3609: coeff = 24'd2226207;
            12'd3610: coeff = 24'd2217482;
            12'd3611: coeff = 24'd2208771;
            12'd3612: coeff = 24'd2200074;
            12'd3613: coeff = 24'd2191392;
            12'd3614: coeff = 24'd2182725;
            12'd3615: coeff = 24'd2174072;
            12'd3616: coeff = 24'd2165434;
            12'd3617: coeff = 24'd2156810;
            12'd3618: coeff = 24'd2148202;
            12'd3619: coeff = 24'd2139608;
            12'd3620: coeff = 24'd2131028;
            12'd3621: coeff = 24'd2122464;
            12'd3622: coeff = 24'd2113914;
            12'd3623: coeff = 24'd2105379;
            12'd3624: coeff = 24'd2096858;
            12'd3625: coeff = 24'd2088353;
            12'd3626: coeff = 24'd2079862;
            12'd3627: coeff = 24'd2071386;
            12'd3628: coeff = 24'd2062925;
            12'd3629: coeff = 24'd2054479;
            12'd3630: coeff = 24'd2046048;
            12'd3631: coeff = 24'd2037632;
            12'd3632: coeff = 24'd2029230;
            12'd3633: coeff = 24'd2020844;
            12'd3634: coeff = 24'd2012473;
            12'd3635: coeff = 24'd2004117;
            12'd3636: coeff = 24'd1995775;
            12'd3637: coeff = 24'd1987449;
            12'd3638: coeff = 24'd1979138;
            12'd3639: coeff = 24'd1970842;
            12'd3640: coeff = 24'd1962561;
            12'd3641: coeff = 24'd1954295;
            12'd3642: coeff = 24'd1946044;
            12'd3643: coeff = 24'd1937809;
            12'd3644: coeff = 24'd1929589;
            12'd3645: coeff = 24'd1921384;
            12'd3646: coeff = 24'd1913194;
            12'd3647: coeff = 24'd1905019;
            12'd3648: coeff = 24'd1896860;
            12'd3649: coeff = 24'd1888716;
            12'd3650: coeff = 24'd1880587;
            12'd3651: coeff = 24'd1872473;
            12'd3652: coeff = 24'd1864375;
            12'd3653: coeff = 24'd1856292;
            12'd3654: coeff = 24'd1848225;
            12'd3655: coeff = 24'd1840173;
            12'd3656: coeff = 24'd1832136;
            12'd3657: coeff = 24'd1824115;
            12'd3658: coeff = 24'd1816110;
            12'd3659: coeff = 24'd1808119;
            12'd3660: coeff = 24'd1800145;
            12'd3661: coeff = 24'd1792185;
            12'd3662: coeff = 24'd1784242;
            12'd3663: coeff = 24'd1776314;
            12'd3664: coeff = 24'd1768401;
            12'd3665: coeff = 24'd1760504;
            12'd3666: coeff = 24'd1752623;
            12'd3667: coeff = 24'd1744757;
            12'd3668: coeff = 24'd1736907;
            12'd3669: coeff = 24'd1729072;
            12'd3670: coeff = 24'd1721254;
            12'd3671: coeff = 24'd1713451;
            12'd3672: coeff = 24'd1705663;
            12'd3673: coeff = 24'd1697892;
            12'd3674: coeff = 24'd1690136;
            12'd3675: coeff = 24'd1682396;
            12'd3676: coeff = 24'd1674671;
            12'd3677: coeff = 24'd1666963;
            12'd3678: coeff = 24'd1659270;
            12'd3679: coeff = 24'd1651593;
            12'd3680: coeff = 24'd1643932;
            12'd3681: coeff = 24'd1636287;
            12'd3682: coeff = 24'd1628658;
            12'd3683: coeff = 24'd1621045;
            12'd3684: coeff = 24'd1613447;
            12'd3685: coeff = 24'd1605866;
            12'd3686: coeff = 24'd1598300;
            12'd3687: coeff = 24'd1590751;
            12'd3688: coeff = 24'd1583217;
            12'd3689: coeff = 24'd1575700;
            12'd3690: coeff = 24'd1568199;
            12'd3691: coeff = 24'd1560713;
            12'd3692: coeff = 24'd1553244;
            12'd3693: coeff = 24'd1545791;
            12'd3694: coeff = 24'd1538354;
            12'd3695: coeff = 24'd1530933;
            12'd3696: coeff = 24'd1523528;
            12'd3697: coeff = 24'd1516139;
            12'd3698: coeff = 24'd1508767;
            12'd3699: coeff = 24'd1501411;
            12'd3700: coeff = 24'd1494071;
            12'd3701: coeff = 24'd1486747;
            12'd3702: coeff = 24'd1479439;
            12'd3703: coeff = 24'd1472148;
            12'd3704: coeff = 24'd1464873;
            12'd3705: coeff = 24'd1457614;
            12'd3706: coeff = 24'd1450372;
            12'd3707: coeff = 24'd1443146;
            12'd3708: coeff = 24'd1435936;
            12'd3709: coeff = 24'd1428743;
            12'd3710: coeff = 24'd1421566;
            12'd3711: coeff = 24'd1414405;
            12'd3712: coeff = 24'd1407261;
            12'd3713: coeff = 24'd1400133;
            12'd3714: coeff = 24'd1393022;
            12'd3715: coeff = 24'd1385927;
            12'd3716: coeff = 24'd1378849;
            12'd3717: coeff = 24'd1371787;
            12'd3718: coeff = 24'd1364742;
            12'd3719: coeff = 24'd1357713;
            12'd3720: coeff = 24'd1350701;
            12'd3721: coeff = 24'd1343706;
            12'd3722: coeff = 24'd1336727;
            12'd3723: coeff = 24'd1329764;
            12'd3724: coeff = 24'd1322818;
            12'd3725: coeff = 24'd1315889;
            12'd3726: coeff = 24'd1308977;
            12'd3727: coeff = 24'd1302081;
            12'd3728: coeff = 24'd1295202;
            12'd3729: coeff = 24'd1288339;
            12'd3730: coeff = 24'd1281493;
            12'd3731: coeff = 24'd1274664;
            12'd3732: coeff = 24'd1267852;
            12'd3733: coeff = 24'd1261057;
            12'd3734: coeff = 24'd1254278;
            12'd3735: coeff = 24'd1247516;
            12'd3736: coeff = 24'd1240771;
            12'd3737: coeff = 24'd1234043;
            12'd3738: coeff = 24'd1227331;
            12'd3739: coeff = 24'd1220637;
            12'd3740: coeff = 24'd1213959;
            12'd3741: coeff = 24'd1207298;
            12'd3742: coeff = 24'd1200654;
            12'd3743: coeff = 24'd1194027;
            12'd3744: coeff = 24'd1187417;
            12'd3745: coeff = 24'd1180824;
            12'd3746: coeff = 24'd1174248;
            12'd3747: coeff = 24'd1167689;
            12'd3748: coeff = 24'd1161147;
            12'd3749: coeff = 24'd1154621;
            12'd3750: coeff = 24'd1148113;
            12'd3751: coeff = 24'd1141622;
            12'd3752: coeff = 24'd1135148;
            12'd3753: coeff = 24'd1128691;
            12'd3754: coeff = 24'd1122252;
            12'd3755: coeff = 24'd1115829;
            12'd3756: coeff = 24'd1109423;
            12'd3757: coeff = 24'd1103035;
            12'd3758: coeff = 24'd1096663;
            12'd3759: coeff = 24'd1090309;
            12'd3760: coeff = 24'd1083972;
            12'd3761: coeff = 24'd1077653;
            12'd3762: coeff = 24'd1071350;
            12'd3763: coeff = 24'd1065065;
            12'd3764: coeff = 24'd1058797;
            12'd3765: coeff = 24'd1052546;
            12'd3766: coeff = 24'd1046312;
            12'd3767: coeff = 24'd1040096;
            12'd3768: coeff = 24'd1033897;
            12'd3769: coeff = 24'd1027715;
            12'd3770: coeff = 24'd1021551;
            12'd3771: coeff = 24'd1015404;
            12'd3772: coeff = 24'd1009274;
            12'd3773: coeff = 24'd1003162;
            12'd3774: coeff = 24'd997067;
            12'd3775: coeff = 24'd990990;
            12'd3776: coeff = 24'd984930;
            12'd3777: coeff = 24'd978887;
            12'd3778: coeff = 24'd972862;
            12'd3779: coeff = 24'd966854;
            12'd3780: coeff = 24'd960864;
            12'd3781: coeff = 24'd954891;
            12'd3782: coeff = 24'd948936;
            12'd3783: coeff = 24'd942998;
            12'd3784: coeff = 24'd937078;
            12'd3785: coeff = 24'd931175;
            12'd3786: coeff = 24'd925290;
            12'd3787: coeff = 24'd919423;
            12'd3788: coeff = 24'd913573;
            12'd3789: coeff = 24'd907740;
            12'd3790: coeff = 24'd901926;
            12'd3791: coeff = 24'd896129;
            12'd3792: coeff = 24'd890349;
            12'd3793: coeff = 24'd884587;
            12'd3794: coeff = 24'd878843;
            12'd3795: coeff = 24'd873117;
            12'd3796: coeff = 24'd867408;
            12'd3797: coeff = 24'd861717;
            12'd3798: coeff = 24'd856043;
            12'd3799: coeff = 24'd850388;
            12'd3800: coeff = 24'd844750;
            12'd3801: coeff = 24'd839130;
            12'd3802: coeff = 24'd833527;
            12'd3803: coeff = 24'd827943;
            12'd3804: coeff = 24'd822376;
            12'd3805: coeff = 24'd816827;
            12'd3806: coeff = 24'd811296;
            12'd3807: coeff = 24'd805783;
            12'd3808: coeff = 24'd800287;
            12'd3809: coeff = 24'd794810;
            12'd3810: coeff = 24'd789350;
            12'd3811: coeff = 24'd783908;
            12'd3812: coeff = 24'd778484;
            12'd3813: coeff = 24'd773078;
            12'd3814: coeff = 24'd767690;
            12'd3815: coeff = 24'd762320;
            12'd3816: coeff = 24'd756968;
            12'd3817: coeff = 24'd751634;
            12'd3818: coeff = 24'd746318;
            12'd3819: coeff = 24'd741019;
            12'd3820: coeff = 24'd735739;
            12'd3821: coeff = 24'd730477;
            12'd3822: coeff = 24'd725233;
            12'd3823: coeff = 24'd720007;
            12'd3824: coeff = 24'd714799;
            12'd3825: coeff = 24'd709609;
            12'd3826: coeff = 24'd704437;
            12'd3827: coeff = 24'd699283;
            12'd3828: coeff = 24'd694147;
            12'd3829: coeff = 24'd689029;
            12'd3830: coeff = 24'd683930;
            12'd3831: coeff = 24'd678849;
            12'd3832: coeff = 24'd673785;
            12'd3833: coeff = 24'd668740;
            12'd3834: coeff = 24'd663713;
            12'd3835: coeff = 24'd658705;
            12'd3836: coeff = 24'd653714;
            12'd3837: coeff = 24'd648742;
            12'd3838: coeff = 24'd643788;
            12'd3839: coeff = 24'd638852;
            12'd3840: coeff = 24'd633935;
            12'd3841: coeff = 24'd629035;
            12'd3842: coeff = 24'd624154;
            12'd3843: coeff = 24'd619291;
            12'd3844: coeff = 24'd614447;
            12'd3845: coeff = 24'd609621;
            12'd3846: coeff = 24'd604813;
            12'd3847: coeff = 24'd600023;
            12'd3848: coeff = 24'd595252;
            12'd3849: coeff = 24'd590499;
            12'd3850: coeff = 24'd585765;
            12'd3851: coeff = 24'd581049;
            12'd3852: coeff = 24'd576351;
            12'd3853: coeff = 24'd571672;
            12'd3854: coeff = 24'd567011;
            12'd3855: coeff = 24'd562368;
            12'd3856: coeff = 24'd557744;
            12'd3857: coeff = 24'd553138;
            12'd3858: coeff = 24'd548551;
            12'd3859: coeff = 24'd543982;
            12'd3860: coeff = 24'd539432;
            12'd3861: coeff = 24'd534900;
            12'd3862: coeff = 24'd530387;
            12'd3863: coeff = 24'd525892;
            12'd3864: coeff = 24'd521416;
            12'd3865: coeff = 24'd516958;
            12'd3866: coeff = 24'd512519;
            12'd3867: coeff = 24'd508098;
            12'd3868: coeff = 24'd503696;
            12'd3869: coeff = 24'd499312;
            12'd3870: coeff = 24'd494947;
            12'd3871: coeff = 24'd490601;
            12'd3872: coeff = 24'd486273;
            12'd3873: coeff = 24'd481963;
            12'd3874: coeff = 24'd477673;
            12'd3875: coeff = 24'd473401;
            12'd3876: coeff = 24'd469147;
            12'd3877: coeff = 24'd464913;
            12'd3878: coeff = 24'd460697;
            12'd3879: coeff = 24'd456499;
            12'd3880: coeff = 24'd452320;
            12'd3881: coeff = 24'd448160;
            12'd3882: coeff = 24'd444019;
            12'd3883: coeff = 24'd439896;
            12'd3884: coeff = 24'd435792;
            12'd3885: coeff = 24'd431707;
            12'd3886: coeff = 24'd427641;
            12'd3887: coeff = 24'd423593;
            12'd3888: coeff = 24'd419564;
            12'd3889: coeff = 24'd415554;
            12'd3890: coeff = 24'd411562;
            12'd3891: coeff = 24'd407589;
            12'd3892: coeff = 24'd403636;
            12'd3893: coeff = 24'd399700;
            12'd3894: coeff = 24'd395784;
            12'd3895: coeff = 24'd391887;
            12'd3896: coeff = 24'd388008;
            12'd3897: coeff = 24'd384148;
            12'd3898: coeff = 24'd380307;
            12'd3899: coeff = 24'd376485;
            12'd3900: coeff = 24'd372682;
            12'd3901: coeff = 24'd368897;
            12'd3902: coeff = 24'd365132;
            12'd3903: coeff = 24'd361385;
            12'd3904: coeff = 24'd357658;
            12'd3905: coeff = 24'd353949;
            12'd3906: coeff = 24'd350259;
            12'd3907: coeff = 24'd346588;
            12'd3908: coeff = 24'd342936;
            12'd3909: coeff = 24'd339303;
            12'd3910: coeff = 24'd335689;
            12'd3911: coeff = 24'd332093;
            12'd3912: coeff = 24'd328517;
            12'd3913: coeff = 24'd324960;
            12'd3914: coeff = 24'd321422;
            12'd3915: coeff = 24'd317902;
            12'd3916: coeff = 24'd314402;
            12'd3917: coeff = 24'd310921;
            12'd3918: coeff = 24'd307459;
            12'd3919: coeff = 24'd304015;
            12'd3920: coeff = 24'd300591;
            12'd3921: coeff = 24'd297186;
            12'd3922: coeff = 24'd293800;
            12'd3923: coeff = 24'd290433;
            12'd3924: coeff = 24'd287085;
            12'd3925: coeff = 24'd283756;
            12'd3926: coeff = 24'd280446;
            12'd3927: coeff = 24'd277156;
            12'd3928: coeff = 24'd273884;
            12'd3929: coeff = 24'd270631;
            12'd3930: coeff = 24'd267398;
            12'd3931: coeff = 24'd264184;
            12'd3932: coeff = 24'd260988;
            12'd3933: coeff = 24'd257812;
            12'd3934: coeff = 24'd254655;
            12'd3935: coeff = 24'd251518;
            12'd3936: coeff = 24'd248399;
            12'd3937: coeff = 24'd245300;
            12'd3938: coeff = 24'd242219;
            12'd3939: coeff = 24'd239158;
            12'd3940: coeff = 24'd236117;
            12'd3941: coeff = 24'd233094;
            12'd3942: coeff = 24'd230090;
            12'd3943: coeff = 24'd227106;
            12'd3944: coeff = 24'd224141;
            12'd3945: coeff = 24'd221195;
            12'd3946: coeff = 24'd218268;
            12'd3947: coeff = 24'd215361;
            12'd3948: coeff = 24'd212473;
            12'd3949: coeff = 24'd209604;
            12'd3950: coeff = 24'd206754;
            12'd3951: coeff = 24'd203924;
            12'd3952: coeff = 24'd201113;
            12'd3953: coeff = 24'd198321;
            12'd3954: coeff = 24'd195548;
            12'd3955: coeff = 24'd192795;
            12'd3956: coeff = 24'd190061;
            12'd3957: coeff = 24'd187347;
            12'd3958: coeff = 24'd184651;
            12'd3959: coeff = 24'd181975;
            12'd3960: coeff = 24'd179318;
            12'd3961: coeff = 24'd176681;
            12'd3962: coeff = 24'd174063;
            12'd3963: coeff = 24'd171464;
            12'd3964: coeff = 24'd168885;
            12'd3965: coeff = 24'd166325;
            12'd3966: coeff = 24'd163784;
            12'd3967: coeff = 24'd161263;
            12'd3968: coeff = 24'd158761;
            12'd3969: coeff = 24'd156278;
            12'd3970: coeff = 24'd153815;
            12'd3971: coeff = 24'd151371;
            12'd3972: coeff = 24'd148947;
            12'd3973: coeff = 24'd146542;
            12'd3974: coeff = 24'd144156;
            12'd3975: coeff = 24'd141790;
            12'd3976: coeff = 24'd139443;
            12'd3977: coeff = 24'd137116;
            12'd3978: coeff = 24'd134808;
            12'd3979: coeff = 24'd132519;
            12'd3980: coeff = 24'd130250;
            12'd3981: coeff = 24'd128001;
            12'd3982: coeff = 24'd125770;
            12'd3983: coeff = 24'd123560;
            12'd3984: coeff = 24'd121368;
            12'd3985: coeff = 24'd119197;
            12'd3986: coeff = 24'd117044;
            12'd3987: coeff = 24'd114911;
            12'd3988: coeff = 24'd112798;
            12'd3989: coeff = 24'd110704;
            12'd3990: coeff = 24'd108630;
            12'd3991: coeff = 24'd106575;
            12'd3992: coeff = 24'd104539;
            12'd3993: coeff = 24'd102523;
            12'd3994: coeff = 24'd100527;
            12'd3995: coeff = 24'd98550;
            12'd3996: coeff = 24'd96593;
            12'd3997: coeff = 24'd94655;
            12'd3998: coeff = 24'd92737;
            12'd3999: coeff = 24'd90838;
            12'd4000: coeff = 24'd88959;
            12'd4001: coeff = 24'd87099;
            12'd4002: coeff = 24'd85259;
            12'd4003: coeff = 24'd83438;
            12'd4004: coeff = 24'd81637;
            12'd4005: coeff = 24'd79855;
            12'd4006: coeff = 24'd78093;
            12'd4007: coeff = 24'd76351;
            12'd4008: coeff = 24'd74628;
            12'd4009: coeff = 24'd72925;
            12'd4010: coeff = 24'd71241;
            12'd4011: coeff = 24'd69577;
            12'd4012: coeff = 24'd67933;
            12'd4013: coeff = 24'd66308;
            12'd4014: coeff = 24'd64702;
            12'd4015: coeff = 24'd63117;
            12'd4016: coeff = 24'd61550;
            12'd4017: coeff = 24'd60004;
            12'd4018: coeff = 24'd58477;
            12'd4019: coeff = 24'd56970;
            12'd4020: coeff = 24'd55482;
            12'd4021: coeff = 24'd54014;
            12'd4022: coeff = 24'd52565;
            12'd4023: coeff = 24'd51136;
            12'd4024: coeff = 24'd49727;
            12'd4025: coeff = 24'd48338;
            12'd4026: coeff = 24'd46968;
            12'd4027: coeff = 24'd45617;
            12'd4028: coeff = 24'd44287;
            12'd4029: coeff = 24'd42976;
            12'd4030: coeff = 24'd41684;
            12'd4031: coeff = 24'd40413;
            12'd4032: coeff = 24'd39161;
            12'd4033: coeff = 24'd37928;
            12'd4034: coeff = 24'd36715;
            12'd4035: coeff = 24'd35522;
            12'd4036: coeff = 24'd34349;
            12'd4037: coeff = 24'd33195;
            12'd4038: coeff = 24'd32061;
            12'd4039: coeff = 24'd30947;
            12'd4040: coeff = 24'd29852;
            12'd4041: coeff = 24'd28777;
            12'd4042: coeff = 24'd27721;
            12'd4043: coeff = 24'd26686;
            12'd4044: coeff = 24'd25670;
            12'd4045: coeff = 24'd24673;
            12'd4046: coeff = 24'd23697;
            12'd4047: coeff = 24'd22740;
            12'd4048: coeff = 24'd21803;
            12'd4049: coeff = 24'd20885;
            12'd4050: coeff = 24'd19987;
            12'd4051: coeff = 24'd19109;
            12'd4052: coeff = 24'd18251;
            12'd4053: coeff = 24'd17412;
            12'd4054: coeff = 24'd16593;
            12'd4055: coeff = 24'd15794;
            12'd4056: coeff = 24'd15014;
            12'd4057: coeff = 24'd14254;
            12'd4058: coeff = 24'd13514;
            12'd4059: coeff = 24'd12794;
            12'd4060: coeff = 24'd12093;
            12'd4061: coeff = 24'd11412;
            12'd4062: coeff = 24'd10750;
            12'd4063: coeff = 24'd10109;
            12'd4064: coeff = 24'd9487;
            12'd4065: coeff = 24'd8885;
            12'd4066: coeff = 24'd8303;
            12'd4067: coeff = 24'd7740;
            12'd4068: coeff = 24'd7197;
            12'd4069: coeff = 24'd6674;
            12'd4070: coeff = 24'd6170;
            12'd4071: coeff = 24'd5687;
            12'd4072: coeff = 24'd5223;
            12'd4073: coeff = 24'd4778;
            12'd4074: coeff = 24'd4354;
            12'd4075: coeff = 24'd3949;
            12'd4076: coeff = 24'd3564;
            12'd4077: coeff = 24'd3199;
            12'd4078: coeff = 24'd2853;
            12'd4079: coeff = 24'd2527;
            12'd4080: coeff = 24'd2221;
            12'd4081: coeff = 24'd1935;
            12'd4082: coeff = 24'd1668;
            12'd4083: coeff = 24'd1421;
            12'd4084: coeff = 24'd1194;
            12'd4085: coeff = 24'd987;
            12'd4086: coeff = 24'd799;
            12'd4087: coeff = 24'd631;
            12'd4088: coeff = 24'd483;
            12'd4089: coeff = 24'd355;
            12'd4090: coeff = 24'd246;
            12'd4091: coeff = 24'd157;
            12'd4092: coeff = 24'd88;
            12'd4093: coeff = 24'd39;
            12'd4094: coeff = 24'd9;
            12'd4095: coeff = 24'd0;
        endcase
    end
endmodule
